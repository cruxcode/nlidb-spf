�� sr -edu.cornell.cs.nlp.spf.parser.ccg.model.Model�5B��B�~ L featureSetst Ljava/util/List;L independentLexicalFeatureSetsq ~ L invalidFeaturest Ljava/util/Set;L lexicont -Ledu/cornell/cs/nlp/spf/ccg/lexicon/ILexicon;L thetat 4Ledu/cornell/cs/nlp/spf/base/hashvector/IHashVector;xpsr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.LinkedList)S]J`�"  xpw   sr Pedu.cornell.cs.nlp.spf.parser.ccg.factoredlex.features.FactoredLexicalFeatureSet�g�պ��� D 
entryScaleI lexemeNextIdD lexemeScaleI nonFactoredNextIdI templateNextIdD templateScaleL entryInitialScorert :Ledu/cornell/cs/nlp/utils/collections/ISerializableScorer;L 	lexemeIdst 5Lit/unimi/dsi/fastutil/objects/Object2IntOpenHashMap;L lexemeInitialScorerq ~ L nonFactoredIdsq ~ L templateIdsq ~ L templateInitialScorerq ~ xr Iedu.cornell.cs.nlp.spf.parser.ccg.model.lexical.AbstractLexicalFeatureSetZ���n3�� Z computeSyntaxAttributeFeaturesL 
featureTagt Ljava/lang/String;L ignoreFiltert Ljava/util/function/Predicate;xp t FACLEXsr !java.lang.invoke.SerializedLambdaoaД,)6� 
I implMethodKind[ capturedArgst [Ljava/lang/Object;L capturingClasst Ljava/lang/Class;L functionalInterfaceClassq ~ L functionalInterfaceMethodNameq ~ L "functionalInterfaceMethodSignatureq ~ L 	implClassq ~ L implMethodNameq ~ L implMethodSignatureq ~ L instantiatedMethodTypeq ~ xp   ur [Ljava.lang.Object;��X�s)l  xp    vr 0edu.cornell.cs.nlp.utils.function.PredicateUtils           xpt java/util/function/Predicatet testt (Ljava/lang/Object;)Zt 0edu/cornell/cs/nlp/utils/function/PredicateUtilst lambda$alwaysTrue$bcad8f2c$1q ~ q ~ ?�         �?�             o?�������sr Eedu.cornell.cs.nlp.spf.parser.ccg.features.basic.scorer.UniformScorerQ�B���S D scorexp        sr 3it.unimi.dsi.fastutil.objects.Object2IntOpenHashMap         F fI sizexr 3it.unimi.dsi.fastutil.objects.AbstractObject2IntMap�o��K<z  xr 8it.unimi.dsi.fastutil.objects.AbstractObject2IntFunction�o��K<z I defRetValuexp    ?@     �sr 9edu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.Lexeme	I����� I hashCodeCacheL 
attributesq ~ L 	constantsq ~ L 
propertiest Ljava/util/Map;L 	signaturet GLedu/cornell/cs/nlp/spf/ccg/lexicon/factored/lambda/FactoringSignature;L tokenst ,Ledu/cornell/cs/nlp/spf/base/token/TokenSeq;xp|��qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sr 0edu.cornell.cs.nlp.spf.mr.lambda.LogicalConstant=Q��� L baseNameq ~ L nameq ~ xr %edu.cornell.cs.nlp.spf.mr.lambda.Term�(G^� L typet .Ledu/cornell/cs/nlp/spf/mr/language/type/Type;xr 2edu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression
n�tL�h  xpsr 3edu.cornell.cs.nlp.spf.mr.language.type.ComplexType� �g��V L domainq ~ 2L rangeq ~ 2xr ,edu.cornell.cs.nlp.spf.mr.language.type.Typeg���� I hashCodeCacheL nameq ~ xp���Nt 
<c,c_pkey>sr 0edu.cornell.cs.nlp.spf.mr.language.type.TermType��6��ǭ L parentt 2Ledu/cornell/cs/nlp/spf/mr/language/type/TermType;xq ~ 6   ct csq ~ 9  �t losq ~ 9   et epsq ~ 9�_Kt c_pkeysq ~ 9 4��t pkeyq ~ ?t pkey_retrievert pkey_retriever:<c,c_pkey>xq ~ /q ~ .sr %java.util.Collections$UnmodifiableMap��t�B L mq ~ (xpsq ~ Gsr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t origint fixed_domainxsr Eedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoringSignature�ڝ�U鞉 I hashCodeI numAttributesL typesq ~ xp|!<    sq ~ sr java.util.ArrayListx����a� I sizexp   w   sq ~ 5|\t <e,e>q ~ ?q ~ ?xq ~ Rsr *edu.cornell.cs.nlp.spf.base.token.TokenSeq�py��An I hashCode[ tokenst [Ljava/lang/String;xp*��ur [Ljava.lang.String;��V��{G  xp   t dehradunw   Fsq ~ '  �Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ _q ~ ^sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~ esq ~ U  uq ~ X   t ofw   Tsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ mq ~ lsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~ ssq ~ U�,Kuq ~ X   t witht thew   sq ~ '�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5"��nt 
<s,s_pkey>sq ~ 9   st sq ~ =sq ~ 9ɬ�;t s_pkeyq ~ Cq ~ Et pkey_retriever:<s,s_pkey>sq ~ 0q ~ �t maharashtrat maharashtra:sxq ~ |q ~ {sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~ �sq ~ U�� puq ~ X   q ~ �w   �sq ~ ';�Чsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~ �sq ~ U;I�uq ~ X   q ~ �t statew   Psq ~ '�F��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t jaipurt jaipur:cxq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~ �sq ~ U�j�uq ~ X   q ~ �w   �sq ~ ' 8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~ �sq ~ U ��uq ~ X   q ~ ww   'sq ~ '\�m�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t 
aurangabadt aurangabad:cxq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~ �sq ~ Ub+$�uq ~ X   q ~ �w   osq ~ '�+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t bhusawalt 
bhusawal:cxq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~ �sq ~ U䲃uq ~ X   q ~ �w   �sq ~ 'h�t'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~ �sq ~ U���uq ~ X   t gurgaonw   sq ~ ' �sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~ �sq ~ U ��uq ~ X   t howw    sq ~ 'k��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5^��pt <<e,t>,<<e,i>,e>>sq ~ 5|-t <e,t>q ~ ?sq ~ 9   tt tpsq ~ 5H��	t 	<<e,i>,e>sq ~ 5|�t <e,i>q ~ ?sq ~ 9   it iq ~ ?q ~ ?t argmaxt argmax:<<e,t>,<<e,i>,e>>xq ~ �q ~ �sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   sq ~ 5W�i�t <<e,t>,<<e,e>,e>>q ~ �sq ~ 5HgKt 	<<e,e>,e>q ~ Sq ~ ?xq ~sq ~ U��uq ~ X   t largestw   Qsq ~ ' 1�Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~"sq ~ U 1�	uq ~ X   t int feetw   7sq ~ '�^��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t kotat kota:cxq ~+q ~*sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~4sq ~ U 2Suq ~ X   q ~-w   �sq ~ '�"l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0sq ~ 5l��t <lo,i>q ~ =q ~t 	elevationt elevation:<lo,i>xq ~;q ~:sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~Fsq ~ U6�0�uq ~ X   t highestw   zsq ~ 'R	+{q ~(sq ~ sq ~ sq ~ 
w   q ~ 4xq ~Mq ~Lsq ~ Gq ~0sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Qq ~5w   sq ~ '�f�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }sq ~ 0q ~ �t haryanat 	haryana:sxq ~Vq ~Usq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~_sq ~ U)�uq ~ X   q ~Xw   �sq ~ '�Ӌ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t 	rishikesht rishikesh:cxq ~fq ~esq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~osq ~ U�F
uq ~ X   q ~hw   �sq ~ 'n��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~vq ~usq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~|sq ~ U 3;�uq ~ X   t mostw   8sq ~ '1�̫sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t katnit katni:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U�Wuq ~ X   q ~�w   isq ~ 'R�}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t deoghart 	deoghar:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~ U\�2uq ~ X   q ~�w   lsq ~ '��]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��t <t,t>q ~q ~t nott 	not:<t,t>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~�sq ~ U  �uq ~ X   t now   Ssq ~ '�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5I:�t 	<<e,t>,i>q ~ �q ~t countt count:<<e,t>,i>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   sq ~ 5I:��t 	<<e,t>,e>q ~ �q ~ ?xq ~�sq ~ U�Xۇuq ~ X   t numberw   Jsq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~=t sizet size:<lo,i>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ U��uq ~ X   q ~w   sq ~ '�I�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t kurukshetrat kurukshetra:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~ UG륏uq ~ X   q ~�w   �sq ~ 'o.F-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ U�q�uq ~ X   q ~ wq ~ �w   6sq ~ '���ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�!��t <b_pkey,<s_pkey,t>>sq ~ 9��-�t b_pkeyq ~ Csq ~ 5I�x�t 
<s_pkey,t>q ~ �q ~t next_tot next_to:<b_pkey,<s_pkey,t>>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N?z��    sq ~ sq ~ Q   w   sq ~ 5?z�t 	<e,<e,t>>q ~ ?q ~ �xq ~sq ~ U���@uq ~ X   t statesw   Ksq ~ '��P�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t argmint argmin:<<e,t>,<<e,i>,e>>xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~sq ~ U!N�uq ~ X   t leastw   ;sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~#q ~"sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~)sq ~ U z�uq ~ X   t arew   sq ~ ' dx.sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~1q ~0sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~7sq ~ U c��uq ~ X   q ~ �t manyw   sq ~ 'POr�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5^��tt <<e,t>,<<e,i>,i>>q ~ �sq ~ 5H���t 	<<e,i>,i>q ~q ~t sumt sum:<<e,t>,<<e,i>,i>>xq ~?q ~>sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~Lsq ~ U�~�Cuq ~ X   t combinedw   3sq ~ 'wr�+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t mumbait mumbai:cxq ~Tq ~Ssq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~]sq ~ U��cuq ~ X   q ~Vw   �sq ~ 'd��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~q ~<xq ~dq ~csq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~jsq ~ U��5�uq ~ X   t lowestw   nsq ~ '�R��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t khandwat 	khandwa:cxq ~rq ~qsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~{sq ~ U�=3�uq ~ X   q ~tw   �sq ~ 'z�G+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t kanpurt kanpur:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U�!&suq ~ X   q ~�w   |sq ~ '��usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ Uk��	uq ~ X   t 	jharkhandw   4sq ~ '�*�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�7��t 	<i,<i,t>>q ~sq ~ 5}�t <i,t>q ~q ~t >t >:<i,<i,t>>q ~<xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N�W9J    sq ~ sq ~ Q   w   q ~	q ~ Sxq ~�sq ~ U6ǁ�uq ~ X   t highert thanw   �sq ~ '��h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t uttar_pradesht uttar_pradesh:sxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~ U�)�uq ~ X   t uttart pradeshw   �sq ~ '�8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�sq ~ UW��uq ~ X   q ~ wq ~w   psq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t jodhpurt 	jodhpur:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~ U�p�"uq ~ X   q ~�w   Rsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ U|ܥuq ~ X   t 
chandigarhw   sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~�sq ~ U��uq ~ X   q ~w   �sq ~ 'ڧXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t reewat reewa:cxq ~ q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~	sq ~ Uu�uq ~ X   q ~w   �sq ~ '�Acsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t nainitalt 
nainital:cxq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~sq ~ Ugj(�uq ~ X   q ~w   vsq ~ '��&sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~ q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~&sq ~ U�C�uq ~ X   t tellt mew   +sq ~ '��}�q ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~.q ~-sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~2q ~�w   sq ~ 'B��?q ~ssq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~6q ~5sq ~ Gq ~xsq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~:q ~}w   �sq ~ '�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~?q ~>sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~Esq ~ U�8muq ~ X   t atq ~t onew   [sq ~ '�Gv�q ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~Mq ~Lsq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Qq ~�w   sq ~ 'A�;�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��}�t <s_pkey,<b_pkey,t>>q ~ �sq ~ 5q�t 
<b_pkey,t>q ~�q ~q ~t next_to:<s_pkey,<b_pkey,t>>xq ~Vq ~Usq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~bsq ~ U��tjuq ~ X   t borderw   �sq ~ 'a���q ~ �sq ~ sq ~ sq ~ 
w   q ~ 4xq ~iq ~hsq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~mq ~ �w   5sq ~ '�.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Wxq ~rq ~qsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~xsq ~ U�b_�uq ~ X   q ~ wq ~ �q ~ hq ~Xw   �sq ~ 'e��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t luckhnowt 
luckhnow:cxq ~q ~~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U�<��uq ~ X   q ~�w   �sq ~ ' /��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U /"�uq ~ X   t doesw   sq ~ 'CG�+q ~ �sq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;q ~ �t 	gurgaon:cxq ~�q ~�sq ~ Gq ~ �sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~ �w   �sq ~ '��$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�sq ~ U��7,uq ~ X   t fewestw   ysq ~ '���ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��t <b_pkey,<t,s_pkey>>q ~�sq ~ 5���ot 
<t,s_pkey>q ~q ~ �q ~t next_to:<b_pkey,<t,s_pkey>>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N@M�4    sq ~ sq ~ Q   w   sq ~ 5@M�Tt 	<e,<t,e>>q ~ ?sq ~ 5���t <t,e>q ~q ~ ?xq ~�sq ~ U���@uq ~ X   q ~w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~ U��]uq ~ X   t smallestw   sq ~ 'b�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t 	darbhangat darbhanga:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U��� uq ~ X   q ~�w   �sq ~ 'B��q ~�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~�t jharkhand:sxq ~�q ~�sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~�w   ssq ~ '@H�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t bhopalt bhopal:cxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U�(�Puq ~ X   q ~�w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~
sq ~ U �uq ~ X   q ~�w   :sq ~ '��Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t 	mussooriet mussoorie:cxq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~sq ~ U)duq ~ X   q ~w   \sq ~ 'E�d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4q ~ �xq ~!q ~ sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~'sq ~ Ubau�uq ~ X   q ~ wq ~ �w   �sq ~ 'OG�q ~<sq ~ sq ~ sq ~ 
w   q ~�xq ~-q ~,sq ~ Gq ~Asq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~1q ~Fw   sq ~ '�}8.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~6q ~5sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~<sq ~ U��5�uq ~ X   q ~mw   _sq ~ '��!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }xq ~Cq ~Bsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Isq ~ U�M0uq ~ X   t biharw   sq ~ '���q ~sq ~ sq ~ sq ~ 
w   q ~ 4q ~xq ~Pq ~Osq ~ Gq ~sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~Tq ~w   �sq ~ '�,�Xq ~Ssq ~ sq ~ sq ~ 
w   q ~Wxq ~Xq ~Wsq ~ Gq ~[sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~\q ~`w   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t jalgaont 	jalgaon:cxq ~aq ~`sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~jsq ~ U���uq ~ X   q ~cw   �sq ~ 'WS�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~pq ~osq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~tq ~�w   esq ~ '��J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Uxq ~yq ~xsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~sq ~ U0�q5uq ~ X   t cityt namedq ~Vw   �sq ~ '�7�q ~sq ~ sq ~ sq ~ 
w   q ~ 4q ~xq ~�q ~�sq ~ Gq ~sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~w   ~sq ~ 'i�Euq ~�sq ~ sq ~ sq ~ 
w   q ~<xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~�w   sq ~ '%���q ~<sq ~ sq ~ sq ~ 
w   q ~�q ~�sq ~ 0q ~t 0t 0:ixq ~�q ~�sq ~ Gq ~Asq ~ N)���    sq ~ sq ~ Q   w   q ~	q ~�q ~ ?xq ~�q ~Fw   �sq ~ 'n�vq ~csq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~ksq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~pw   sq ~ '2�^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~=t 
populationt population:<lo,i>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ U�b�uq ~ X   q ~�w   Nsq ~ '�Ղ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~�sq ~ U 3�uq ~ X   t doq ~�w   ksq ~ '����q ~sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~�w   �sq ~ '�|۸q ~Qsq ~ sq ~ sq ~ 
w   q ~Uxq ~�q ~�sq ~ Gq ~Ysq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~^w   �sq ~ 'B��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~�sq ~ U i�uq ~ X   q ~ wq ~w   wsq ~ '��,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }sq ~ 0q ~ �t madhya_pradesht madhya_pradesh:sxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U�uuq ~ X   t madhyaq ~�w   �sq ~ 'A�r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~ Uz�p�uq ~ X   t sparsestw   Osq ~ '�hНsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5^-֟t <b_pkey,s_pkey>q ~�q ~ �q ~t next_to:<b_pkey,s_pkey>xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~ U��tjuq ~ X   q ~ew   sq ~ 'nw4q ~@sq ~ sq ~ sq ~ 
w   q ~ }sq ~ 0q ~ �q ~Lt bihar:sxq ~q ~sq ~ Gq ~Esq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~q ~Jw   �sq ~ 'W��q ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~q ~sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~#q ~�w   Gsq ~ '�Jz�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~(q ~'sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~.sq ~ U i�uq ~ X   q ~ wq ~w   �sq ~ '3>
�q ~@sq ~ sq ~ sq ~ 
w   q ~xq ~4q ~3sq ~ Gq ~Esq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~8q ~Jw   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~q ~�xq ~=q ~<sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~Csq ~ U!N�uq ~ X   q ~w   asq ~ 'Z#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~Jq ~Isq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Psq ~ U�<��uq ~ X   t nagpurw   sq ~ ' 19�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~Xq ~Wsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~^sq ~ U 0��uq ~ X   t havew   sq ~ '�D�zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~fq ~esq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~lsq ~ U c��uq ~ X   q ~ �q ~:w   ^sq ~ '�i8q ~(sq ~ sq ~ sq ~ 
w   q ~,xq ~rq ~qsq ~ Gq ~0sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~vq ~5w   �sq ~ 'ȼ��q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~zq ~ysq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~~q ~�w   �sq ~ '�@�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U�@(uq ~ X   t pleasew   sq ~ '�Ӭxq ~^sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~fsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~kw   sq ~ '���q ~sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~�w   (sq ~ '��nQq ~�sq ~ sq ~ sq ~ 
w   q ~<q ~<xq ~�q ~�sq ~ Gq ~�sq ~ No��    sq ~ sq ~ Q   w   q ~ Sq ~ Sxq ~�q ~�w   �sq ~ '�5�6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~ UW��uq ~ X   q ~ wq ~w   Wsq ~ '��I�q ~vsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~{sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~�w   
sq ~ 'ǥ\q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~�q ~�w   Dsq ~ '�AXq ~sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~w   sq ~ 'xq ~ ,sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;q ~ Zt 
dehradun:cxq ~�q ~�sq ~ Gq ~ Isq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~ Ww   �sq ~ '�<2q ~:sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~?sq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�q ~Dw   xsq ~ '�3� q ~�sq ~ sq ~ sq ~ 
w   q ~ }q ~�xq ~�q ~�sq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~�w   �sq ~ ',�?�q ~<sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~�q ~�sq ~ Gq ~Asq ~ N�ǂ    sq ~ sq ~ Q   w   q ~	q ~�xq ~�q ~Fw   �sq ~ '�C�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ U�0��uq ~ X   t 	rajasthanw   sq ~ '�<�kq ~ �sq ~ sq ~ sq ~ 
w   q ~ 4q ~ �xq ~�q ~�sq ~ Gq ~ �sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~q ~ �w   �sq ~ '�8N[q ~sq ~ sq ~ sq ~ 
w   q ~ 4xq ~q ~sq ~ Gq ~#sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	q ~(w   	sq ~ '�Ԝxq ~�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;q ~�t chandigarh:cxq ~q ~sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~q ~�w   Csq ~ 'H�'8q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~q ~�w   �sq ~ '���q ~vsq ~ sq ~ sq ~ 
w   q ~ 4q ~Uxq ~q ~sq ~ Gq ~{sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~#q ~�w   �sq ~ '��[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~(q ~'sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~.sq ~ U��tjuq ~ X   q ~ew   Usq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~5q ~4sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~;sq ~ U6�0�uq ~ X   q ~Iw   Zsq ~ '��
q ~ �sq ~ sq ~ sq ~ 
w   q ~ 4xq ~Aq ~@sq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Eq ~ �w   !sq ~ 'QHܹq ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~Iq ~Hsq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~Mq ~�w   ]sq ~ 'PG�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;t patnat patna:cxq ~Rq ~Qsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~[sq ~ UX!�uq ~ X   q ~Tw   usq ~ 'X.�@q ~Osq ~ sq ~ sq ~ 
w   q ~ 4xq ~aq ~`sq ~ Gq ~Wsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~eq ~\w   sq ~ ' 8)Csq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~jq ~isq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~psq ~ U 7�uq ~ X   q ~ vw   Lsq ~ '{ɡq ~�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~�t rajasthan:sxq ~vq ~usq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~|q ~�w   �sq ~ 'ȆB�q ~ ysq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~sq ~ Gq ~ �sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~ �w   csq ~ '+u4)q ~osq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gq ~tsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~yw   %sq ~ '  x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U   �uq ~ X   t aw   }sq ~ 'c�5Nq ~�sq ~ sq ~ sq ~ 
w   q ~�q ~<q ~<xq ~�q ~�sq ~ Gq ~�sq ~ N���    sq ~ sq ~ Q   w   q ~	q ~ Sq ~ Sxq ~�q ~�w   �sq ~ 'XLÆq ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~
w   -sq ~ '%Nq ~osq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~wsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~|w   sq ~ 'П�~q ~Ssq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gq ~[sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~`w   1sq ~ '�^�8q ~Gsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;q ~St nagpur:cxq ~�q ~�sq ~ Gq ~Lsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~Qw   �sq ~ 'i���q ~8sq ~ sq ~ sq ~ 
w   q ~<xq ~�q ~�sq ~ Gq ~Bsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~Gw   sq ~ 'g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~ U�+X�uq ~ X   t biggestw   &sq ~ 'Ü��q ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~xq ~�q ~�sq ~ Gq ~sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~
w   Asq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~ U��cuq ~ X   t ranchiw   *sq ~ '\�)q ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Gq ~#sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~(w   �sq ~ 'z��q ~Qsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~Ysq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~ q ~^w   )sq ~ ' 8#Asq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~sq ~ U 7�uq ~ X   t whatw   sq ~ '��n�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�sq ~ 0q ~	t equalst equals:<e,<e,t>>xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N�Uܘ    sq ~ sq ~ Q   w   q ~�q ~	xq ~sq ~ Ud��Uuq ~ X   t 	excludingw   �sq ~ ':�-+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4sq ~ 0q ~ ;t noidat noida:cxq ~$q ~#sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~-sq ~ UB%�uq ~ X   q ~&w   �sq ~ '�ʋq ~�sq ~ sq ~ sq ~ 
w   q ~ }q ~wxq ~3q ~2sq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~7q ~�w   rsq ~ 'ZR<�q ~ �sq ~ sq ~ sq ~ 
w   q ~�xq ~;q ~:sq ~ Gq ~ �sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~?q ~ �w   fsq ~ '�Q��q ~<sq ~ sq ~ sq ~ 
w   q ~�xq ~Cq ~Bsq ~ Gq ~Asq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~Gq ~Fw   �sq ~ '~9kq ~�sq ~ sq ~ sq ~ 
w   q ~ }q ~�xq ~Kq ~Jsq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~Oq ~�w   �sq ~ '�\�Xq ~osq ~ sq ~ sq ~ 
w   q ~sxq ~Sq ~Rsq ~ Gq ~wsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~Wq ~|w   �sq ~ 'V��q ~<sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~[q ~Zsq ~ Gq ~Asq ~ N���    sq ~ sq ~ Q   w   q ~�q ~ ?xq ~_q ~Fw   �sq ~ '��\q ~�sq ~ sq ~ sq ~ 
w   q ~ }q ~ �xq ~cq ~bsq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~gq ~�w   �sq ~ ':�l�q ~sq ~ sq ~ sq ~ 
w   q ~xq ~kq ~jsq ~ Gq ~sq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~oq ~w   tsq ~ '��w�q ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~sq ~rsq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~wq ~�w   "sq ~ 'w#�q ~ �sq ~ sq ~ sq ~ 
w   q ~ }q ~ �xq ~{q ~zsq ~ Gq ~ �sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~q ~ �w   �sq ~ 'b�q ~�sq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~�w   >sq ~ 'n���q ~ ysq ~ sq ~ sq ~ 
w   q ~ }xq ~�q ~�sq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~ �w   dsq ~ '��A�q ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~xq ~�q ~�sq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~�w   �sq ~ 'x�J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~�sq ~ U��]uq ~ X   q ~�w   �sq ~ '���q ~asq ~ sq ~ sq ~ 
w   q ~<xq ~�q ~�sq ~ Gq ~fsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~kw   9sq ~ '�Cdq ~�sq ~ sq ~ sq ~ 
w   q ~q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~�q ~�w   �sq ~ '���q ~�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ;q ~�t ranchi:cxq ~�q ~�sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~�w   �sq ~ 'n�B�q ~%sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Gq ~*sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�q ~/w   2sq ~ '�B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U��[uq ~ X   t whichw   $sq ~ 'ڿt�q ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~�xq ~�q ~�sq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~�w   �sq ~ '@�eq ~ �sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~ �w   sq ~ '�?��q ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~�xq ~�q ~�sq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~�w   �sq ~ 'cٔ�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~�w    sq ~ '��ژsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~�sq ~ U��7,uq ~ X   q ~�w   �sq ~ '� ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~sq ~ U  huq ~ X   t isw   Bsq ~ '��g�q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~q ~sq ~ Gq ~ �sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~q ~ �w   bsq ~ '&pxq ~|sq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~q ~�w   �sq ~ '9=�q ~Osq ~ sq ~ sq ~ 
w   q ~ 4q ~Sxq ~#q ~"sq ~ Gq ~Wsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~'q ~\w   hsq ~ 'Q���q ~!sq ~ sq ~ sq ~ 
w   q ~%xq ~+q ~*sq ~ Gq ~)sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~/q ~.w   jsq ~ 'I �q ~<sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~3q ~2sq ~ Gq ~Asq ~ N��S    sq ~ sq ~ Q   w   q ~	q ~ ?xq ~7q ~Fw   Ysq ~ 'ؖE�q ~ ,sq ~ sq ~ sq ~ 
w   q ~ 4q ~�xq ~;q ~:sq ~ Gq ~ Isq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~?q ~ Ww   �sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~Dq ~Csq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~Jsq ~ U  huq ~ X   q ~w   sq ~ 'eIq ~|sq ~ sq ~ sq ~ 
w   q ~ 4xq ~Pq ~Osq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Tq ~�w   0sq ~ 'y�Ƙq ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~Xq ~Wsq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~\q ~�w   �sq ~ '�l
�q ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~`q ~_sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~dq ~�w   .sq ~ '�TP�q ~Gsq ~ sq ~ sq ~ 
w   q ~ 4q ~�xq ~hq ~gsq ~ Gq ~Lsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~lq ~Qw   �sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~qq ~psq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~wsq ~ U  �uq ~ X   t byw   #sq ~ ';Wvq ~osq ~ sq ~ sq ~ 
w   q ~ }q ~Wxq ~~q ~}sq ~ Gq ~tsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�q ~yw   �sq ~ 'OS;\q ~sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~sq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~�q ~w   gsq ~ ' 6Szsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U 5�;uq ~ X   t showw   Esq ~ '�>͜sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~t truet true:txq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  T    sq ~ sq ~ Q   w   q ~xq ~�sq ~ U�Jpuq ~ X   q ~,t therew   �sq ~ ' 6�$sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U 6M�uq ~ X   t thatw   qsq ~ '�݋sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ }sq ~ 0q ~ �t 
uttrakhandt uttrakhand:sxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~�sq ~ U �_tuq ~ X   q ~�w   Xsq ~ '��q ~^sq ~ sq ~ sq ~ 
w   q ~bxq ~�q ~�sq ~ Gq ~fsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~kw   Vsq ~ '�˴q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~�w   �sq ~ 'Ԍӌq ~�sq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�q ~�w   sq ~ '��٤sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~ U��aeuq ~ X   q ~%t metersw   sq ~ '���Xq ~csq ~ sq ~ sq ~ 
w   q ~gxq ~�q ~�sq ~ Gq ~ksq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�q ~pw   `sq ~ 'z�9jq ~�sq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Gq ~�sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�q ~ w   @sq ~ '�\��q ~ �sq ~ sq ~ sq ~ 
w   q ~ }xq ~	q ~	 sq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	q ~ �w   /sq ~ 'E�Kq ~ �sq ~ sq ~ sq ~ 
w   q ~ 4q ~ �xq ~		q ~	sq ~ Gq ~ �sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~	q ~ �w   �sq ~ 'X��q ~!sq ~ sq ~ sq ~ 
w   q ~ 4xq ~	q ~	sq ~ Gq ~)sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	q ~.w   ?sq ~ 'z���q ~sq ~ sq ~ sq ~ 
w   q ~ 4xq ~	q ~	sq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	q ~w   ,sq ~ '��3�q ~�sq ~ sq ~ sq ~ 
w   q ~ }xq ~	!q ~	 sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	%q ~�w   Hsq ~ ' 0�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~	*q ~	)sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~	0sq ~ U 0R/uq ~ X   t cant youw   Msq ~ '}��+q ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~�xq ~	8q ~	7sq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~	<q ~�w   =sq ~ '{g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@xq ~	Aq ~	@sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~	Gsq ~ U�ۂuq ~ X   t totalw   <sq ~ ';�#Kq ~�sq ~ sq ~ sq ~ 
w   q ~ 4q ~�xq ~	Nq ~	Msq ~ Gq ~�sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~	Rq ~�w   {sq ~ '���q ~�sq ~ sq ~ sq ~ 
w   q ~ }xq ~	Vq ~	Usq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	Zq ~�w   Isq ~ '�)Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	_q ~	^sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~	esq ~ U 3;�uq ~ X   q ~w   mxsq ~ !        sq ~ #    ?@      xsq ~ #    ?@     osr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.LexicalTemplateg��%��	 I hashCodeL 	argumentsq ~ L 
propertiesq ~ (L 	signatureq ~ )L templatet 0Ledu/cornell/cs/nlp/spf/ccg/categories/Category;xpYY�Qsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t #0<<e,t>,e>t #0<<e,t>,e>:<<e,t>,e>xq ~	pq ~	osq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~	ysr 5edu.cornell.cs.nlp.spf.ccg.categories.ComplexCategory�f�Ք�nl I hashCodeCacheL syntaxt <Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/ComplexSyntax;xr .edu.cornell.cs.nlp.spf.ccg.categories.CategorycK=�.A� L 	semanticst Ljava/lang/Object;xpsr 'edu.cornell.cs.nlp.spf.mr.lambda.Lambda��Kβ�� L argumentt +Ledu/cornell/cs/nlp/spf/mr/lambda/Variable;L bodyt 4Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L typet 5Ledu/cornell/cs/nlp/spf/mr/language/type/ComplexType;xq ~ 3sr )edu.cornell.cs.nlp.spf.mr.lambda.Variable�u#$rP L 	singletonq ~ xq ~ 1q ~ �sr 5it.unimi.dsi.fastutil.objects.ReferenceSets$Singleton�7y�J| L elementq ~	}xpq ~	�sq ~	sq ~	�q ~ �sq ~	�q ~	�sr (edu.cornell.cs.nlp.spf.mr.lambda.Literalŕtb��� [ 	argumentst 5[Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L 	predicateq ~	�[ 	signaturet /[Ledu/cornell/cs/nlp/spf/mr/language/type/Type;L typeq ~ 2xq ~ 3ur 5[Ledu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression;|�㰢�[i  xp   sq ~	sq ~	�q ~ ?sq ~	�q ~	�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~	�sr ;it.unimi.dsi.fastutil.objects.ReferenceSets$UnmodifiableSet�7y�J|  xr Iit.unimi.dsi.fastutil.objects.ReferenceCollections$UnmodifiableCollection�7y�J| L 
collectiont 3Lit/unimi/dsi/fastutil/objects/ReferenceCollection;xpsr 2it.unimi.dsi.fastutil.objects.ReferenceOpenHashSet         F fI sizexp?@     q ~	�q ~	�xq ~	�ur /[Ledu.cornell.cs.nlp.spf.mr.language.type.Type;>L5��  xp   q ~ ?q ~sq ~	�uq ~	�   q ~	�sq ~	�sq ~	�?@     q ~	�q ~	�xq ~	�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~	�q ~	�q ~	�xsq ~ 0sr <edu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType&��M
� I minArgsZ orderSensitiveL optiont ELedu/cornell/cs/nlp/spf/mr/language/type/RecursiveComplexType$Option;xq ~ 5l�6�t <t*,t>q ~q ~    sr Cedu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType$Option�^g� �� Z isOrderSensitiveI 
minNumArgsxp    t andt 
and:<t*,t>uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~	�q ~	�xq ~ �q ~	�q ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~	�xq ~�sr 4it.unimi.dsi.fastutil.objects.ReferenceSets$EmptySet�7y�J|  xpsq ~ 5q~Et <<e,t>,<<e,t>,e>>q ~ �q ~�n�]sr :edu.cornell.cs.nlp.spf.ccg.categories.syntax.ComplexSyntax$���q\P^ I hashCodeI 	numSlahesL leftt 5Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax;L rightq ~	�L slasht 4Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Slash;xr 3edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntaxʊ�	�|��  xp8���   sq ~	��k�   sr @edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntax$SimpleSyntax��eBg� I hashCodeL 	attributeq ~ L labelq ~ xq ~	� 3�t nonet Ssq ~	�ȠU�   q ~	�sq ~	� 4�wq ~	�t NPsr 2edu.cornell.cs.nlp.spf.ccg.categories.syntax.Slashѕ�����> C cxp \sq ~	� /sq ~	� 3�kq ~	�t Nq ~	�w   Gsq ~	k{r�|sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ St #0<e,e>t #0<e,e>:<e,e>xq ~	�q ~	�sq ~ Gq ~Ysq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	�sr 4edu.cornell.cs.nlp.spf.ccg.categories.SimpleCategory��4_C� I hashCodeCacheL syntaxt BLedu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax$SimpleSyntax;xq ~	|sq ~	�uq ~	�   q ~Uq ~	�q ~	�uq ~	�   q ~ ?q ~ ?4m�Pq ~	�w   sq ~	kS	 {sq ~ sq ~ sq ~ 
w   q ~	�xq ~	�q ~	�sq ~ Gq ~wsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	�sq ~	�sq ~	�uq ~	�   q ~sq ~	�q ~	�uq ~	�   q ~ ?q ~ ?GOq ~	�w   Asq ~	k�Yޣsq ~ sq ~ sq ~ 
w   q ~	�xq ~	�q ~	�sq ~ Gq ~ksq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	�sq ~	�sq ~	�uq ~	�   q ~gq ~	�q ~	�uq ~	�   q ~ ?q ~ ?�Uwq ~	�w   sq ~	k�RVpsq ~ sq ~ sq ~ 
w   q ~	�xq ~	�q ~	�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~	�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?VM}Dq ~	�w   sq ~	k�m��sq ~ sq ~ sq ~ 
w   q ~	�xq ~
q ~
sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~
sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?�h��q ~	�w   sq ~	k~W�sq ~ sq ~ sq ~ 
w    xq ~
q ~
sq ~ Gq ~Fsq ~ N  �    sq ~ sq ~ Q    w    xq ~
sq ~	zsq ~	sq ~	�q ~�sq ~	�q ~
sq ~	sq ~	�q ~ �sq ~	�q ~
sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~
sq ~	�uq ~	�   q ~
sq ~	�sq ~	�?@     q ~
q ~
xq ~
uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~
xq ~ �sq ~	�sq ~	�?@     q ~
q ~
xq ~
uq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~
xq ~�q ~	�sq ~ 5�~t <<<e,t>,e>,<<e,t>,e>>q ~�q ~�~W�!sq ~	����z   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	��ƥY   q ~	�q ~	�q ~	�q ~	�w   sq ~	kYE�sq ~ sq ~ sq ~ 
w   q ~	qxq ~
5q ~
4sq ~ Gq ~hsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~
9sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~
<sq ~	sq ~	�q ~ �sq ~	�q ~
?sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~
Dsq ~	�uq ~	�   sq ~	�uq ~	�   q ~
Dsq ~	�sq ~	�?@     q ~
<q ~
Dxq ~
<uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~
Dsq ~	�sq ~	�?@     q ~
?q ~
Dxq ~
?uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~
?q ~
<q ~
Dxq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~
?q ~
<xq ~ �q ~
Uq ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~
<xq ~�q ~	�q ~	�nu
�sq ~	�8���   sq ~	��f   q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   ]sq ~	k~0�sq ~ sq ~ sq ~ 
w   q ~	�xq ~
`q ~
_sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~
dsq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?7+?�q ~	�w   sq ~	k,���sq ~ sq ~ sq ~ 
w    xq ~
lq ~
ksq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~
rsq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~
usq ~	sq ~	�q ~ ?sq ~	�q ~
xsq ~	�uq ~	�   q ~
xsq ~	�sq ~	�?@     q ~
uq ~
xxq ~
uuq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~
uxq ~ �q ~	�sq ~ 5JW`Lt <<e,t>,<e,t>>q ~ �q ~ �,���sq ~	��9�   sq ~	� 4��q ~	�t PPq ~
�q ~	�w   ,sq ~	k<��sq ~ sq ~ sq ~ 
w   q ~	�sq ~ 0q ~ St #1<e,e>t #1<e,e>:<e,e>xq ~
�q ~
�sq ~ Gq ~�sq ~ No��    sq ~ sq ~ Q   w   q ~ Sq ~ Sxq ~
�sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~
�sq ~	sq ~	�q ~ ?sq ~	�q ~
�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~
�q ~
�q ~	�uq ~	�   q ~ ?q ~ ?sq ~	�uq ~	�   q ~
�q ~
�q ~
�uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	BEsq ~	��P�   q ~
�q ~	�q ~	�w   gsq ~	kV�$�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~t #0<<e,t>,<<e,e>,e>>t %#0<<e,t>,<<e,e>,e>>:<<e,t>,<<e,e>,e>>xq ~
�q ~
�sq ~ Gq ~fsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~
�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~
�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~
�sq ~	�uq ~	�   q ~
�sq ~	�sq ~	�?@     q ~
�q ~
�xq ~
�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~
�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~<uq ~	�   q ~ =q ~q ~	�q ~q ~
�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?q ~	�q ~��j�sq ~	��ƥY   q ~	�q ~	�q ~	�w   ;sq ~	k 	��sq ~ sq ~ sq ~ 
w   q ~
�xq ~
�q ~
�sq ~ Gq ~�sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~
�sq ~	zsq ~	sq ~	�q ~sq ~	�q ~
�sq ~	sq ~	�q ~ �sq ~	�q ~
�sq ~	sq ~	�q ~ �sq ~	�q ~
�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~
�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~
�sq ~	�sq ~	�?@     q ~
�q ~
�xq ~
�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~
�sq ~	�sq ~	�?@     q ~
�q ~
�xq ~
�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~
�q ~
�q ~
�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~
�q ~
�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~�uq ~	�   q ~ =q ~q ~	�q ~q ~
�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~
�xq ~�q ~	�q ~	�sq ~	�sq ~	�?@      xsq ~ 5˹�)t <<e,i>,<<e,t>,<<e,t>,e>>>q ~q ~	����Esq ~	��]�   sq ~	��ƥY   q ~	�q ~	�q ~	�q ~
�q ~	�w   5sq ~	kI�Ssq ~ sq ~ sq ~ 
w   q ~
�xq ~q ~sq ~ Gq ~sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~
sq ~	sq ~	�q ~ Ssq ~	�q ~sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~
q ~xq ~
uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~
xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~q ~xq ~uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~xq ~ Ssq ~	�sq ~	�?@     q ~
q ~xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~
xq ~q ~	�q ~�a�sq ~	�����   sq ~	��ƥY   q ~	�q ~	�q ~	�q ~	�q ~	�w   Tsq ~	k�;�sq ~ sq ~ sq ~ 
w    xq ~/q ~.sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~5sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~8sq ~	sq ~	�q ~ �sq ~	�q ~;sq ~	sq ~	�q ~ ?sq ~	�q ~>sq ~	�uq ~	�   sq ~	�uq ~	�   q ~>sq ~	�sq ~	�?@     q ~>q ~8xq ~8uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~>sq ~	�sq ~	�?@     q ~>q ~;xq ~;uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~>q ~8q ~;xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~8q ~;xq ~ �sq ~	�sq ~	�?@     q ~8xq ~
�q ~	�sq ~ 5˪xt <<e,t>,<<e,t>,<e,t>>>q ~ �q ~
��;�%sq ~	�8���   sq ~	��f   q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   Fsq ~	ks�sq ~ sq ~ sq ~ 
w   q ~	�xq ~[q ~Zsq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~_sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~bsq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~gsq ~	�uq ~	�   q ~gsq ~	�sq ~	�?@     q ~gq ~bxq ~buq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~bxq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~qsq ~	�uq ~	�   q ~qq ~rq ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~nq ~ �uq ~	�   q ~ �q ~q ~ ?q ~	�q ~��n��sq ~	��ƥY   q ~	�q ~	�q ~	�w   sq ~	k����sq ~ sq ~ sq ~ 
w   q ~	�xq ~{q ~zsq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~	�sq ~	�uq ~	�   q ~q ~	�q ~	�uq ~	�   q ~ ?q ~ ?���q ~	�w   
sq ~	k���sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~sq ~	�q ~�q ~�q ~	�q ~����sq ~	��|��   q ~	�q ~	�q ~	�w   2sq ~	k�	�@sq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t #0<t,t>t #0<t,t>:<t,t>sq ~ 0q ~	t #0<e,<e,t>>t #0<e,<e,t>>:<e,<e,t>>xq ~�q ~�sq ~ Gq ~sq ~ N�Uܘ    sq ~ sq ~ Q   w   q ~�q ~	xq ~�sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?q ~q ~�q ~�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~	_p�sq ~	��P�   q ~
�q ~	�q ~	�w   csq ~	k����sq ~ sq ~ sq ~ 
w   q ~
�q ~	�xq ~�q ~�sq ~ Gq ~fsq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~�sq ~	zsq ~	q ~
�sq ~	�uq ~	�   q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~
�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?q ~	�q ~�Z`O�q ~
�w   bsq ~	k�գ�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~
��՟�sq ~	�mLߍ   sq ~	�ȠU�   q ~	�q ~	�q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�w   Msq ~	k��sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?��|q ~	�w   (sq ~	kW��sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?zǋq ~	�w   -sq ~	k���Ssq ~ sq ~ sq ~ 
w   q ~	qxq ~�q ~�sq ~ Gq ~�sq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~sq ~	sq ~	�q ~	sq ~	�q ~sq ~	sq ~	�q ~ �sq ~	�q ~sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~q ~xq ~uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~q ~xq ~uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~q ~q ~xq ~uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~q ~q ~xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~q ~q ~xq ~ �q ~,q ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~q ~xq ~ Ssq ~	�sq ~	�?@     q ~q ~q ~xq ~ �uq ~	�   q ~ �q ~q ~ ?sq ~	�sq ~	�?@     q ~q ~xq ~�sq ~	�sq ~	�?@     q ~xsq ~ 5�Ї�t <<e,<e,t>>,<<e,t>,e>>q ~	q ~�q ~	�sq ~ 5{�t <<e,t>,<<e,<e,t>>,<<e,t>,e>>>q ~ �q ~8�
�_sq ~	��<�   sq ~	���;!   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	�(Iɟ   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   ^sq ~	k�L(�sq ~ sq ~ sq ~ 
w   q ~	�xq ~Dq ~Csq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Hsq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~<uq ~	�   q ~ =q ~sq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	�GOaq ~
�w   #sq ~	kx�sq ~ sq ~ sq ~ 
w    xq ~Yq ~Xsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~_sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~bsq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~gsq ~	�uq ~	�   q ~gsq ~	�sq ~	�?@     q ~bq ~gxq ~buq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~bxq ~ �q ~nsq ~ 0q ~�q ~ wt the:<<e,t>,e>uq ~	�   q ~ �q ~ ?q ~	�q ~�x~'sq ~	��ƥY   q ~	�q ~	�q ~	�w   sq ~	kw%�bsq ~ sq ~ sq ~ 
w    xq ~wq ~vsq ~ Gq ~ssq ~ N  �    sq ~ sq ~ Q    w    xq ~{sq ~	zsq ~	sq ~	�q ~ Ssq ~	�q ~~sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~~q ~�xq ~~uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~~xq ~ Sq ~	�sq ~ 5�T��t <<e,e>,<e,e>>q ~ Sq ~ Sw%��sq ~	��z�M   q ~	�q ~	�q ~	�w   4sq ~	kK��"sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~q ~�q ~�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~
���sq ~	��9�   q ~
�q ~
�q ~	�w   Usq ~	kB�V�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ?t #0et #0e:exq ~�q ~�sq ~ Gq ~�sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~ }uq ~	�   q ~ �q ~ �>�:q ~	�w   Hsq ~	k�E�"sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~q ~�q ~�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~
�!d��sq ~	�mLߍ   sq ~	�ȠU�   q ~	�q ~	�q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�w   Vsq ~	k���5sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gq ~sq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~�q ~�q ~	�q ~ S��}Usq ~	��|�   q ~	�q ~	�q ~	�w   Esq ~	k��{@sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~*sq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~�sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~	�9��sq ~	�(Iɟ   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�w   Jsq ~	k��{@sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~sq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~ sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~q ~xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~xq ~ �q ~	�q ~	�9��sq ~	�(Iɟ   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�w   Isq ~	k���sq ~ sq ~ sq ~ 
w   q ~	qxq ~q ~sq ~ Gq ~Asq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~sq ~	sq ~	�q ~	sq ~	�q ~sq ~	sq ~	�q ~ ?sq ~	�q ~!sq ~	�uq ~	�   sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~(sq ~	�uq ~	�   sq ~	�uq ~	�   q ~(sq ~	�sq ~	�?@     q ~(q ~xq ~uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~(q ~!sq ~	�sq ~	�?@     q ~q ~(q ~!xq ~uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~(q ~!q ~xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~!q ~q ~xq ~ �q ~9q ~	quq ~	�   q ~ �q ~ ?q ~�q ~9q ~�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xsq ~ 5���t <<e,<e,t>>,<e,t>>q ~	q ~ �q ~	�sq ~ 5�"(tt <<e,t>,<<e,<e,t>>,<e,t>>>q ~ �q ~A	�i(sq ~	��7F   sq ~	���   sq ~	�ȠU�   q ~	�q ~	�q ~	�sq ~	�(Iɟ   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   Ysq ~	k���sq ~ sq ~ sq ~ 
w   q ~	�xq ~Mq ~Lsq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Qsq ~	�sq ~	�uq ~	�   q ~q ~	�q ~	�uq ~	�   q ~ ?q ~ ?E�֒q ~	�w   sq ~	k�уsq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~Yq ~Xsq ~ Gq ~Asq ~ N��S    sq ~ sq ~ Q   w   q ~	q ~ ?xq ~]sq ~	zsq ~	q ~sq ~	q ~sq ~	q ~!sq ~	�uq ~	�   sq ~	�uq ~	�   q ~'q ~9q ~�uq ~	�   q ~ �q ~q ~�q ~9q ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xq ~Aq ~	�q ~C.r�q ~Ew   Osq ~	k���	sq ~ sq ~ sq ~ 
w   q ~	�xq ~oq ~nsq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~ssq ~	�sq ~	�uq ~	�   q ~ �q ~	�q ~	�uq ~	�   q ~ ?q ~ ?Z���q ~	�w   sq ~	k�d�sq ~ sq ~ sq ~ 
w   q ~	�xq ~{q ~zsq ~ Gq ~Esq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~	�sq ~	�uq ~	�   q ~q ~	�q ~	�uq ~	�   q ~ ?q ~ ?�{��q ~	�w   6sq ~	k(�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gq ~�sq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~
�(�>sq ~	��|��   q ~	�q ~	�q ~	�w   	sq ~	kk�ƹsq ~ sq ~ sq ~ 
w   q ~
�q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~�sq ~	zsq ~	sq ~	�q ~ Ssq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�q ~�q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~�xq ~�q ~	�q ~	�sq ~	�sq ~	�?@      xsq ~ 5�U�%t <<e,e>,<<e,t>,<<e,t>,e>>>q ~ Sq ~	�7!�sq ~	��]�   sq ~	��ƥY   q ~	�q ~	�q ~	�q ~
�q ~	�w   Xsq ~	k����sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~sq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	q ~�sq ~	q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~uq ~	�   q ~ ?q ~ ?q ~q ~�q ~�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~	 ��~q ~�w   7sq ~	k4W��sq ~ sq ~ sq ~ 
w   q ~
�q ~	qxq ~�q ~�sq ~ Gq ~�sq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~	sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~�q ~xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~q ~�q ~xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~�q ~�q ~xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�q ~xq ~ �q ~q ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~ Ssq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~�sq ~	�sq ~	�?@     q ~�xq ~8q ~	�q ~:[�B�sq ~	��<�   sq ~	���;!   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	�(Iɟ   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   Ssq ~	k�2.dsq ~ sq ~ sq ~ 
w   q ~
�xq ~0q ~/sq ~ Gq ~�sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~4sq ~	zsq ~	sq ~	�q ~ Ssq ~	�q ~7sq ~	sq ~	�q ~ �sq ~	�q ~:sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~?sq ~	�uq ~	�   q ~?sq ~	�sq ~	�?@     q ~:q ~?xq ~:uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~:xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~Isq ~	�uq ~	�   q ~Isq ~	�sq ~	�?@     q ~7q ~Ixq ~7uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~7xq ~ Ssq ~	�sq ~	�?@     q ~7q ~:xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~7xq ~�q ~	�sq ~ 5wй�t <<e,e>,<<e,t>,e>>q ~ Sq ~�!���sq ~	�����   sq ~	��ƥY   q ~	�q ~	�q ~	�q ~	�q ~	�w   sq ~	k�h��sq ~ sq ~ sq ~ 
w    xq ~^q ~]sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~dsq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~gq ~gq ~	�q ~ S�h�sq ~	���!�   q ~	�q ~	�q ~	�w   sq ~	k@�H�sq ~ sq ~ sq ~ 
w   q ~�xq ~mq ~lsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~ssq ~	�q ~�9|vq ~	�w   nsq ~	k��sq ~ sq ~ sq ~ 
w   q ~	�xq ~xq ~wsq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~|sq ~	�sq ~	�uq ~	�   q ~wq ~	�q ~	�uq ~	�   q ~ ?q ~ ?t��Yq ~	�w    sq ~	k�
Y�sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~)sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~%q ~	�q ~	�uq ~	�   q ~ ?q ~ ?j�pq ~	�w   .sq ~	k>�#sq ~ sq ~ sq ~ 
w   q ~	qxq ~�q ~�sq ~ Gq ~*sq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~	sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~�q ~�sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�q ~�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~ �q ~�q ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~ Ssq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~ �uq ~	�   q ~ �q ~q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~�sq ~	�sq ~	�?@     q ~�xq ~8q ~	�q ~:SBl/sq ~	�='S   sq ~	��w��   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	��P�   q ~
�q ~	�q ~	�q ~	�q ~	�q ~	�w   Wsq ~	kIJ�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~t #0tt #0t:txq ~�q ~�sq ~ Gq ~�sq ~ N  T    sq ~ sq ~ Q   w   q ~xq ~�sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~�q ~�sq ~	�sq ~	�?@      xq ~ �
��ksq ~	�ȠU�   q ~	�q ~	�q ~	�w   ksq ~	k:��sq ~ sq ~ sq ~ 
w   q ~
�xq ~�q ~�sq ~ Gq ~*sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~	zsq ~	q ~�sq ~	q ~�sq ~	q ~�sq ~	�uq ~	�   q ~�sq ~	q ~�sq ~	�uq ~	�   q ~�q ~�q ~�uq ~	�   q ~ �q ~sq ~	�sq ~	�?@     q ~�q ~�xq ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~�sq ~	�sq ~	�?@     q ~�xq ~8q ~	�q ~:��q ~�w   Rsq ~	kn�g@sq ~ sq ~ sq ~ 
w   q ~	qxq ~q ~sq ~ Gq ~�sq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~	sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~	q ~xq ~	uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~	xq ~ �q ~q ~	quq ~	�   q ~ �q ~ ?q ~	�q ~Ä#�Lsq ~	��|�(   q ~	�q ~	�q ~	�w   Psq ~	k��Ysq ~ sq ~ sq ~ 
w   q ~
�xq ~q ~sq ~ Gq ~�sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~ sq ~	zsq ~	q ~�sq ~	q ~�sq ~	q ~�sq ~	�uq ~	�   q ~�sq ~	q ~�sq ~	�uq ~	�   q ~�q ~�q ~�uq ~	�   q ~ =q ~q ~	�q ~q ~�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~�xq ~�q ~	�q ~	�sq ~	�sq ~	�?@      xq ~΋#R�q ~�w   /sq ~	k�[Bsq ~ sq ~ sq ~ 
w   q ~	�xq ~3q ~2sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~7sq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~
�q ~uq ~	�   q ~ �q ~q ~ ?sq ~	�sq ~	�?@     q ~
�xq ~�q ~	�q ~	�sq ~	�sq ~	�?@      xq ~
�˨�q ~
�w   'sq ~	kp�sq ~ sq ~ sq ~ 
w   q ~	�xq ~Jq ~Isq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Nsq ~	�sq ~	�uq ~	�   q ~ �q ~	�q ~	�uq ~	�   q ~ ?q ~ ?)�7�q ~	�w   sq ~	k�[sq ~ sq ~ sq ~ 
w   q ~	�xq ~Vq ~Usq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Zsq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~]sq ~	�uq ~	�   q ~]q ~^q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ SjVB�sq ~	���!�   q ~	�q ~	�q ~	�w   sq ~	k�K�sq ~ sq ~ sq ~ 
w   q ~�q ~	�q ~
�xq ~fq ~esq ~ Gq ~�sq ~ N���    sq ~ sq ~ Q   w   q ~	q ~ Sq ~ Sxq ~jsq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~
�q ~
�q ~	�uq ~	�   q ~ ?q ~ ?sq ~	�uq ~	�   q ~
�q ~
�q ~
�uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	$��q ~
�w   hsq ~	k��S7sq ~ sq ~ sq ~ 
w   q ~	�xq ~~q ~}sq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~ �q ~	�q ~	�uq ~	�   q ~ ?q ~ ?��zq ~	�w   sq ~	k�ҀQsq ~ sq ~ sq ~ 
w   q ~
�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�q ~�q ~�uq ~	�   q ~ =q ~q ~	�q ~q ~�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?q ~	�q ~�dQ�sq ~	��ƥY   q ~	�q ~	�q ~	�w   Ksq ~	k1�j�sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?����q ~	�w   %sq ~	k���sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�xq ~ �sq ~	�sq ~	�?@     q ~�xq ~
�q ~	�q ~S���sq ~	��g�   sq ~	��z�z   q ~	�q ~	�q ~	�q ~	�q ~	�w   Dsq ~	k��msq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?|	�Aq ~	�w   sq ~	k8/[�sq ~ sq ~ sq ~ 
w   q ~	qxq ~�q ~�sq ~ Gq ~?sq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~	sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~	sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~�q ~xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~q ~	sq ~	�sq ~	�?@     q ~�q ~	q ~xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~	q ~xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~	q ~�q ~�xq ~ �q ~q ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~ Ssq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~uq ~	�   q ~ �q ~q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~�sq ~	�sq ~	�?@     q ~�xq ~8q ~	�q ~:M^�sq ~	�='S   sq ~	��w��   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	��P�   q ~
�q ~	�q ~	�q ~	�q ~	�q ~	�w   Qsq ~	kG�sq ~ sq ~ sq ~ 
w   q ~
�xq ~2q ~1sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~6sq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~
�q ~
�q ~<uq ~	�   q ~ =q ~q ~
�sq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	�h*q ~
�w   sq ~	kq�*�sq ~ sq ~ sq ~ 
w    xq ~Gq ~Fsq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~Msq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~Psq ~	sq ~	�q ~ ?sq ~	�q ~Ssq ~	�uq ~	�   q ~Ssq ~	�sq ~	�?@     q ~Pq ~Sxq ~Puq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~Pxq ~ �q ~	�q ~
�q�'sq ~	�	f�   q ~
�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�w   ?sq ~	kT��!sq ~ sq ~ sq ~ 
w   q ~�xq ~aq ~`sq ~ Gq ~Asq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~esq ~	zsq ~	q ~sq ~	q ~sq ~	q ~!sq ~	�uq ~	�   q ~dq ~�q ~9q ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xq ~Aq ~	�q ~CS�0�q ~Ew   sq ~	k��)sq ~ sq ~ sq ~ 
w   q ~	qq ~�xq ~tq ~ssq ~ Gq ~Asq ~ N���    sq ~ sq ~ Q   w   q ~�q ~ ?xq ~xsq ~	zsq ~	q ~sq ~	q ~sq ~	q ~!sq ~	�uq ~	�   q ~%q ~�q ~9q ~�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xq ~Aq ~	�q ~C��@q ~Ew   lsq ~	k�+9Tsq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	zsq ~	q ~�sq ~	q ~�sq ~	q ~�sq ~	�uq ~	�   q ~�sq ~	q ~�sq ~	�uq ~	�   q ~�q ~�q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~�q ~ �uq ~	�   q ~ �q ~q ~ ?sq ~	�sq ~	�?@     q ~�xq ~�q ~	�q ~	�sq ~	�sq ~	�?@      xq ~Ο&`(q ~�w   3sq ~	k����sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?u��q ~	�w   0sq ~	kjw�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~�sq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~�sq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~<q ~Nsq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	��q ~
�w   Csq ~	k@#{�sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~q ~	�q ~	�uq ~	�   q ~ ?q ~ ?���q ~	�w   sq ~	k���(sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~0sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~,q ~	�q ~	�uq ~	�   q ~ ?q ~ ?m��q ~	�w   $sq ~	kiQsq ~ sq ~ sq ~ 
w   q ~�q ~	qxq ~�q ~�sq ~ Gq ~Asq ~ N�ǂ    sq ~ sq ~ Q   w   q ~	q ~�xq ~�sq ~	zsq ~	q ~sq ~	q ~sq ~	q ~!sq ~	�uq ~	�   q ~%q ~�q ~9q ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xq ~Aq ~	�q ~ChIqq ~Ew   jsq ~	k�P3�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gq ~sq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�xq ~ �sq ~	�sq ~	�?@     q ~�xq ~
�q ~	�q ~S�P/�sq ~	�8���   sq ~	��k�   q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   sq ~	k��o�sq ~ sq ~ sq ~ 
w   q ~	�xq ~q ~sq ~ Gq ~[sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~	�sq ~	�uq ~	�   q ~Wq ~	�q ~	�uq ~	�   q ~ ?q ~ ?@��q ~	�w   =sq ~	k�7�msq ~ sq ~ sq ~ 
w   q ~	�xq ~q ~sq ~ Gq ~Wsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~	�sq ~	�uq ~	�   q ~Sq ~	�q ~	�uq ~	�   q ~ ?q ~ ?;2�Aq ~	�w   :sq ~	k��v�sq ~ sq ~ sq ~ 
w    xq ~'q ~&sq ~ Gq ~%sq ~ N  �    sq ~ sq ~ Q    w    xq ~+sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~.sq ~	sq ~	�q ~ ?sq ~	�q ~1sq ~	�uq ~	�   q ~1sq ~	�sq ~	�?@     q ~.q ~1xq ~.uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~.xq ~ �q ~	�q ~
���r�sq ~	�(J�]   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~
�q ~	�w   &sq ~	kGsJ�sq ~ sq ~ sq ~ 
w   q ~�xq ~?q ~>sq ~ Gq ~sq ~ N���    sq ~ sq ~ Q   w   q ~�xq ~Csq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~Fsq ~	sq ~	�q ~ ?sq ~	�q ~Isq ~	�uq ~	�   sq ~	�uq ~	�   q ~Isq ~	�sq ~	�?@     q ~Iq ~Fxq ~Fuq ~	�   q ~ ?q ~q ~Oq ~�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~Fxq ~ �q ~	�q ~
�|�[�sq ~	��z�M   q ~	�q ~	�q ~	�w   [sq ~	kܞf�sq ~ sq ~ sq ~ 
w   q ~	�xq ~Yq ~Xsq ~ Gq ~ �sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~]sq ~	�sq ~	�uq ~	�   q ~ �q ~	�q ~	�uq ~	�   q ~ ?q ~ ?���pq ~	�w   *sq ~	kf{!sq ~ sq ~ sq ~ 
w   q ~	�xq ~eq ~dsq ~ Gq ~ Isq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~isq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?vG�q ~	�w   9sq ~	kq�%{sq ~ sq ~ sq ~ 
w    xq ~qq ~psq ~ Gq ~�sq ~ N  �    sq ~ sq ~ Q    w    xq ~usq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~xsq ~	sq ~	�q ~ ?sq ~	�q ~{sq ~	�uq ~	�   q ~{sq ~	�sq ~	�?@     q ~{q ~xxq ~xuq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~xxq ~ �q ~	�q ~
�q�!�sq ~	�	aJ   q ~
�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�w   +sq ~	k)U$�sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?�PK�q ~	�w   sq ~	k�y��sq ~ sq ~ sq ~ 
w   q ~
�xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~	zsq ~	sq ~	�q ~ Ssq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~�xq ~ Ssq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~�sq ~	�sq ~	�?@     q ~�xq ~	�q ~	�q ~�\�sq ~	�(��O   sq ~	��]�   sq ~	��ƥY   q ~	�q ~	�q ~	�q ~
�q ~	�q ~	�q ~	�w   8sq ~	k��B�sq ~ sq ~ sq ~ 
w   q ~�q ~	qq ~�xq ~�q ~�sq ~ Gq ~Asq ~ N)���    sq ~ sq ~ Q   w   q ~	q ~�q ~ ?xq ~�sq ~	zsq ~	q ~sq ~	q ~sq ~	q ~!sq ~	�uq ~	�   sq ~	�uq ~	�   q ~'q ~9q ~	quq ~	�   q ~ �q ~ ?q ~�q ~9q ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xq ~Aq ~	�q ~CB��q ~Ew   asq ~	k���^sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~
����~sq ~	�mL1-   sq ~	�ȠU�   q ~	�q ~	�q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�w   !sq ~	kn@��sq ~ sq ~ sq ~ 
w   q ~	�xq ~q ~sq ~ Gq ~sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~	�sq ~	�uq ~	�   q ~q ~	�q ~	�uq ~	�   q ~ ?q ~ ?';�Yq ~	�w   sq ~	k(W~sq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Gq ~ �sq ~ N  �    sq ~ sq ~ Q    w    xq ~sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~q ~xq ~uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~xq ~ �q ~	�q ~
�(S�sq ~	��z�M   q ~	�q ~	�q ~	�w   sq ~	k��2"sq ~ sq ~ sq ~ 
w   q ~	�xq ~'q ~&sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~+sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?U�X�q ~	�w   sq ~	kÏn�sq ~ sq ~ sq ~ 
w   q ~
�q ~	qxq ~3q ~2sq ~ Gq ~xsq ~ N���    sq ~ sq ~ Q   w   q ~q ~�xq ~7sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~:sq ~	sq ~	�q ~	sq ~	�q ~=sq ~	sq ~	�q ~ �sq ~	�q ~@sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~Esq ~	�uq ~	�   q ~Esq ~	�sq ~	�?@     q ~@q ~Exq ~@uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~@xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~Osq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~Tsq ~	�uq ~	�   sq ~	�uq ~	�   q ~Tsq ~	�sq ~	�?@     q ~Tq ~:xq ~:uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~Tq ~Osq ~	�sq ~	�?@     q ~Oq ~Tq ~=xq ~=uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~Oq ~Tq ~=q ~:xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~Oq ~:q ~=xq ~ �q ~eq ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~=q ~:xq ~ Ssq ~	�sq ~	�?@     q ~@q ~=q ~:xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~=q ~:xq ~�sq ~	�sq ~	�?@     q ~:xq ~8q ~	�q ~:�.-�sq ~	�='S   sq ~	��w��   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	��P�   q ~
�q ~	�q ~	�q ~	�q ~	�q ~	�w   \sq ~	kG0�Hsq ~ sq ~ sq ~ 
w   q ~�xq ~xq ~wsq ~ Gq ~sq ~ N?z��    sq ~ sq ~ Q   w   q ~	xq ~|sq ~	zsq ~	q ~�sq ~	q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?q ~q ~�q ~�uq ~	�   q ~q ~sq ~	�sq ~	�?@     q ~�xq ~ �q ~	�q ~	Fx��q ~�w   dsq ~	k�^�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~Asq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~	zsq ~	q ~sq ~	q ~sq ~	q ~!sq ~	�uq ~	�   q ~dq ~�q ~9q ~�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~q ~xq ~ �sq ~	�sq ~	�?@     q ~xq ~Aq ~	�q ~C���|q ~Ew   Bsq ~	k�H��sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~fsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~bq ~	�q ~	�uq ~	�   q ~ ?q ~ ?�C�yq ~	�w   sq ~	k��p�sq ~ sq ~ sq ~ 
w   q ~	qxq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ NI:�t    sq ~ sq ~ Q   w   q ~�xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~	sq ~	�q ~�sq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�uq ~	�   q ~�q ~�sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�q ~�xq ~	�uq ~	�   q ~q ~q ~sq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~ �q ~�q ~	quq ~	�   q ~ �q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~ Ssq ~	�sq ~	�?@     q ~�q ~�q ~�xq ~uq ~	�   q ~ �q ~q ~ ?sq ~	�sq ~	�?@     q ~�q ~�xq ~�sq ~	�sq ~	�?@     q ~�xq ~8q ~	�q ~:�&��sq ~	��<�   sq ~	���;!   sq ~	��ƥ�   q ~	�q ~	�q ~	�sq ~	�(Iɟ   sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�q ~	�w   `sq ~	krS{�sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~Lsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?+N��q ~	�w   )sq ~	kl�b�sq ~ sq ~ sq ~ 
w   q ~	�xq ~ q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?%��`q ~	�w   "sq ~	kʆ�sq ~ sq ~ sq ~ 
w   q ~�q ~	�xq ~q ~sq ~ Gq ~�sq ~ N�W9J    sq ~ sq ~ Q   w   q ~	q ~ Sxq ~sq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�q ~Nsq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	mG��q ~
�w   msq ~	k���sq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N  �    sq ~ sq ~ Q    w    xq ~$sq ~	zsq ~	sq ~	�q ~sq ~	�q ~'q ~'q ~	�q ~����sq ~	��|�   q ~	�q ~	�q ~	�w   @sq ~	k��sq ~ sq ~ sq ~ 
w    xq ~-q ~,sq ~ Gq ~�sq ~ N  �    sq ~ sq ~ Q    w    xq ~1sq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~4q ~4q ~	�q ~ S���sq ~	�ȠU�   q ~	�q ~	�q ~	�w   Zsq ~	k(�Ysq ~ sq ~ sq ~ 
w    xq ~:q ~9sq ~ Gq ~�sq ~ N  �    sq ~ sq ~ Q    w    xq ~>sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~Asq ~	sq ~	�q ~ ?sq ~	�q ~Dsq ~	�uq ~	�   q ~Dsq ~	�sq ~	�?@     q ~Aq ~Dxq ~Auq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~Axq ~ �q ~	�q ~
�(�ysq ~	��|�(   q ~	�q ~	�q ~	�w   sq ~	k�O�sq ~ sq ~ sq ~ 
w   q ~	�xq ~Qq ~Psq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~Usq ~	zsq ~	sq ~	�q ~ ?sq ~	�q ~Xsq ~	�uq ~	�   q ~Xq ~Yq ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sfv�sq ~	�ȠU�   q ~	�q ~	�q ~	�w   sq ~	kȨ�sq ~ sq ~ sq ~ 
w   q ~	�xq ~aq ~`sq ~ Gq ~fsq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~esq ~	zsq ~	q ~
�sq ~	�uq ~	�   q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~
�q ~uq ~	�   q ~ �q ~q ~ ?q ~	�q ~Á�9�q ~
�w   sq ~	k��sq ~ sq ~ sq ~ 
w   q ~	�q ~�xq ~rq ~qsq ~ Gq ~ �sq ~ Nl�    sq ~ sq ~ Q   w   q ~ Sq ~ ?xq ~vsq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?ڄs�q ~	�w   <sq ~	kTB�|sq ~ sq ~ sq ~ 
w   q ~	�xq ~~q ~}sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?=�Pq ~	�w   1sq ~	kI�Gmsq ~ sq ~ sq ~ 
w   q ~
�xq ~�q ~�sq ~ Gq ~Hsq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~�sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~�sq ~	sq ~	�q ~ Ssq ~	�q ~�sq ~	�uq ~	�   sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~�xq ~ �sq ~	sq ~	�q ~ ?sq ~	�q ~�sq ~	�uq ~	�   q ~�sq ~	�sq ~	�?@     q ~�q ~�xq ~�uq ~	�   q ~ ?q ~ ?sq ~	�sq ~	�?@     q ~�xq ~ Ssq ~	�sq ~	�?@     q ~�q ~�xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~�xq ~q ~	�q ~�a��sq ~	�����   sq ~	��ƥ�   q ~	�q ~	�q ~	�q ~	�q ~	�w   Nsq ~	kL�Zsq ~ sq ~ sq ~ 
w   q ~�q ~
�xq ~�q ~�sq ~ Gq ~�sq ~ N�W9J    sq ~ sq ~ Q   w   q ~	q ~ Sxq ~�sq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~<q ~
�sq ~	�sq ~	�?@     q ~
�q ~
�xq ~�uq ~	�   q ~ ?q ~ ?q ~sq ~	�sq ~	�?@     q ~
�xq ~ �q ~	�q ~	Ċ��q ~
�w   esq ~	k�n9sq ~ sq ~ sq ~ 
w   q ~
�q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N�C�j    sq ~ sq ~ Q   w   q ~q ~ Sxq ~�sq ~	zsq ~	q ~
�sq ~	q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�sq ~	q ~
�sq ~	�uq ~	�   q ~
�q ~
�q ~	�uq ~	�   q ~ ?q ~ ?q ~	�q ~ Sq ~
�q ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~
�xq ~�q ~	�q ~	�sq ~	�sq ~	�?@      xq ~
�iw�Aq ~
�w   _sq ~	k�CЭsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Gq ~ �sq ~ N  E    sq ~ sq ~ Q   w   q ~ ?xq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~ 4uq ~	�   q ~ ;q ~ A��Jq ~	�w   Lsq ~	kW��sq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~�sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?�<�q ~	�w   >sq ~	k�̱%sq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t #0<e,<t,e>>t #0<e,<t,e>>:<e,<t,e>>xq ~�q ~�sq ~ Gsq ~ Gsq ~ J?@     w      q ~ Lq ~ Mxsq ~ N@M�4    sq ~ sq ~ Q   w   q ~�xq ~ sq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~sq ~	sq ~	�q ~ ?sq ~	�q ~sq ~	�uq ~	�   q ~sq ~	�uq ~	�   q ~sq ~	�sq ~	�?@     q ~q ~xq ~uq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~q ~xq ~�uq ~	�   q ~ ?q ~q ~ ?sq ~	�sq ~	�?@     q ~xq ~ Sq ~	�sq ~ 5JW'�t <<e,t>,<e,e>>q ~ �q ~ S�K��sq ~	���
�   q ~	�q ~
�q ~	�w   fsq ~	k~��sq ~ sq ~ sq ~ 
w   q ~
�xq ~q ~sq ~ Gq ~�sq ~ NW�m�    sq ~ sq ~ Q   w   q ~xq ~sq ~	zsq ~	q ~sq ~	q ~sq ~	q ~sq ~	�uq ~	�   q ~sq ~	q ~sq ~	�uq ~	�   q ~q ~,q ~�uq ~	�   q ~ �q ~sq ~	�sq ~	�?@     q ~q ~xq ~sq ~	�sq ~	�?@     q ~q ~q ~xq ~
�uq ~	�   q ~ �q ~ Sq ~ ?sq ~	�sq ~	�?@     q ~q ~xq ~�sq ~	�sq ~	�?@     q ~xq ~8q ~	�q ~:�8q ~<w    sq ~	k/�sq ~ sq ~ sq ~ 
w   q ~	�xq ~5q ~4sq ~ Gq ~�sq ~ N|!<    sq ~ sq ~ Q   w   q ~ Sxq ~9sq ~	�sq ~	�uq ~	�   q ~�q ~	�q ~	�uq ~	�   q ~ ?q ~ ?���q ~	�w   sq ~	k��Usq ~ sq ~ sq ~ 
w   q ~�xq ~Aq ~@sq ~ Gq ~�sq ~ N@M�4    sq ~ sq ~ Q   w   q ~�xq ~Esq ~	zsq ~	sq ~	�q ~ �sq ~	�q ~Hsq ~	sq ~	�q ~ ?sq ~	�q ~Ksq ~	�uq ~	�   q ~Ksq ~	�uq ~	�   q ~Ksq ~	�sq ~	�?@     q ~Hq ~Kxq ~Huq ~	�   q ~ ?q ~sq ~	�sq ~	�?@     q ~Hq ~Kxq ~�uq ~	�   q ~ ?q ~q ~ ?sq ~	�sq ~	�?@     q ~Hxq ~ Sq ~	�q ~�N$!sq ~	��7�   q ~	�sq ~	�ȠU�   q ~	�q ~	�q ~	�q ~	�w   ixsq ~ !        sr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCoordinationFeatureSet�4tHWcg+ Z cpapFeaturesZ cpp1FeaturesZ reptFeaturesxpsr Dedu.cornell.cs.nlp.spf.parser.ccg.features.basic.RuleUsageFeatureSet�k�d�L2� D scaleZ unaryRulesOnlyL 	ignoreSetq ~ xp?������� sr java.util.HashSet�D�����4  xpw   ?@      xsr Ledu.cornell.cs.nlp.spf.parser.ccg.features.basic.DynamicWordSkippingFeatures%�q�� L emptyCategoryq ~	lL 
featureTagq ~ xpsq ~	�p    sq ~	�zT�lq ~	�t EMPTYt DYNSKIPxq ~ sq ~ sq ~ Q   w   q ~ xq ~isr %java.util.Collections$UnmodifiableSet��я��U  xq ~ sq ~`w   ?@     sr .edu.cornell.cs.nlp.spf.base.hashvector.KeyArgs���]e.ɘ I hashCodeL arg1q ~ L arg2q ~ L arg3q ~ L arg4q ~ L arg5q ~ xp2Iݬq ~ t 
TMPDEFAULTpppsq ~mwzq ~ t XEMEDEFAULTpppsq ~m'��q ~ t 
LEXDEFAULTpppxsr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoredLexicon�>�"z L lexemesq ~ (L lexemesByTypeq ~ (L 	templatesq ~ (xpsq ~ J?@     `w   �   Tq ~ �sq ~`w   ?@     q ~ �q ~8q ~�xq ~�sq ~`w   ?@     q ~�q ~�q ~�xq ~sq ~`w   ?@     q ~�q ~q ~�xq ~Dsq ~`w   ?@     q ~�q ~9q ~xq ~�sq ~`w   ?@     q ~ �q ~�q ~�xq ~ tsq ~`w   ?@     q ~ ixq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~]q ~�q ~	Kxq ~Qsq ~`w   ?@     q ~Fq ~�q ~exq ~\sq ~`w   ?@     q ~ q ~^q ~Nxq ~msq ~`w   ?@     q ~-q ~bxq ~�sq ~`w   ?@     q ~�q ~�xq ~�sq ~`w   ?@     q ~�xq ~(sq ~`w   ?@     q ~q ~q ~�xq ~ �sq ~`w   ?@     q ~ �xq ~sq ~`w   ?@     q ~ xq ~*sq ~`w   ?@     q ~xq ~ �sq ~`w   ?@     q ~�q ~�q ~ �xq ~	Hsq ~`w   ?@     q ~	=xq ~xsq ~`w   ?@     q ~mxq ~ fsq ~`w   ?@     q ~ [xq ~�sq ~`w   ?@     q ~�q ~Uq ~�xq ~ �sq ~`w   ?@     q ~ xq ~�q ~}xq ~_sq ~`w   ?@     q ~Txq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�xq ~	1sq ~`w   ?@     q ~	&xq ~`sq ~`w   ?@     q ~�q ~Uq ~Rxq ~�sq ~`w   ?@     q ~�q ~Hq ~�xq ~�sq ~`w   ?@     q ~�xq ~Jsq ~`w   ?@     q ~?q ~1q ~xq ~�sq ~`w   ?@     q ~�q ~�q ~�xq ~�sq ~`w   ?@     q ~�q ~�q ~
xq ~ �sq ~`w   ?@     q ~ �xq ~�sq ~`w   ?@     q ~�q ~�q ~�xq ~�sq ~`w   ?@     q ~�xq ~qsq ~`w   ?@     q ~fxq ~ Wsq ~`w   ?@     q ~�q ~ +q ~8xq ~ �sq ~`w   ?@     q ~ �q ~	q ~>xq ~sq ~`w   ?@     q ~xq ~ �sq ~`w   ?@     q ~�q ~xq ~ �xq ~Fsq ~`w   ?@     q ~;q ~Xq ~�q ~�q ~@q ~0q ~*xq ~#sq ~`w   ?@     q ~xq ~psq ~`w   ?@     q ~�q ~bq ~�xq ~Msq ~`w   ?@     q ~;xq ~5sq ~`w   ?@     q ~oq ~Jq ~'xq ~.sq ~`w   ?@     q ~ q ~	q ~(xq ~�sq ~`w   ?@     q ~q ~q ~�xq ~^sq ~`w   ?@     q ~�q ~�q ~Pxq ~�sq ~`w   ?@     q ~�q ~�q ~	xq ~�sq ~`w   ?@     q ~�q ~�q ~Jxq ~�sq ~`w   ?@     q ~�q ~�q ~~xq ~�sq ~`w   ?@     q ~�xq ~sq ~`w   ?@     q ~hq ~q ~�xq ~�sq ~`w   ?@     q ~�q ~�q ~�q ~�q ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�q ~wq ~`xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~sq ~0q ~�xq ~ysq ~`w   ?@     q ~nq ~�q ~{xq ~|sq ~`w   ?@     q ~Pq ~nq ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~q ~Mq ~{xq ~sq ~`w   ?@     q ~Mq ~q ~	xq ~�sq ~`w   ?@     q ~�q ~�q ~+xq ~�sq ~`w   ?@     q ~uq ~q ~�xq ~�sq ~`w   ?@     q ~�xq ~sq ~`w   ?@     q ~q ~Rq ~$xq ~ �sq ~`w   ?@     q ~fq ~q ~ �xq ~�sq ~`w   ?@     q ~xq ~Ksq ~`w   ?@     q ~q ~@xq ~�sq ~`w   ?@     q ~�xq ~
sq ~`w   ?@     q ~�q ~�q ~�xq ~ksq ~`w   ?@     q ~`q ~�q ~2xq ~ksq ~`w   ?@     q ~�q ~]q ~�xq ~�sq ~`w   ?@     q ~�q ~�q ~	5xq ~�sq ~`w   ?@     q ~Fq ~	Sq ~�xq ~}sq ~`w   ?@     q ~rq ~	[q ~3xq ~<sq ~`w   ?@     q ~1q ~�q ~7xq ~'sq ~`w   ?@     q ~xq ~�sq ~`w   ?@     q ~pq ~�q ~mxq ~�sq ~`w   ?@     q ~�q ~�q ~�xq ~/sq ~`w   ?@     q ~$q ~�q ~�xq ~�sq ~`w   ?@     q ~�xxsq ~ J?@     w       q ~8sq ~`w   ?@     q ~�q ~9q ~�q ~�q ~3xq ~�sq ~`w   @?@     .q ~�q ~�q ~�q ~�q ~pq ~�q ~�q ~�q ~Jq ~�q ~�q ~>q ~�q ~	q ~fq ~�q ~�q ~Mq ~�q ~�q ~�q ~q ~�q ~�q ~]q ~�q ~�q ~�q ~q ~^q ~	q ~Fq ~ �q ~Jq ~�q ~q ~?q ~	q ~�q ~�q ~+q ~	Sq ~�q ~ +q ~�q ~�xq ~�sq ~`w   ?@     q ~�xq ~	sq ~`w    ?@     q ~�q ~�q ~@q ~q ~-q ~ iq ~ �q ~�q ~ �q ~q ~�q ~q ~ [q ~mq ~Tq ~q ~q ~�q ~fq ~	&q ~�xq ~ �sq ~`w   @?@     (q ~nq ~Pq ~�q ~�q ~q ~mq ~�q ~(q ~ �q ~�q ~oq ~sq ~�q ~�q ~�q ~wq ~�q ~�q ~�q ~q ~}q ~Nq ~uq ~�q ~�q ~1q ~q ~@q ~8q ~
q ~Fq ~�q ~Uq ~ �q ~q ~Uq ~�q ~q ~ �q ~�xq ~�sq ~`w   ?@     q ~�xq ~5sq ~`w   ?@     q ~0xq ~]sq ~`w   ?@     q ~Xxq ~�sq ~`w   ?@     q ~`q ~�q ~�q ~7xq ~�sq ~`w   @?@     'q ~ q ~�q ~q ~0q ~]q ~{q ~{q ~	Kq ~�q ~�q ~Mq ~�q ~�q ~�q ~bq ~nq ~Pq ~~q ~�q ~q ~ �q ~`q ~	q ~�q ~Rq ~�q ~�q ~ xq ~�q ~'q ~	5q ~ q ~xq ~Hq ~�q ~q ~8q ~eq ~�xq ~sq ~`w   ?@     q ~xq ~/sq ~`w   ?@     q ~hq ~�q ~q ~Rq ~�q ~*q ~$xq ~�sq ~`w   ?@     q ~�q ~;q ~�q ~$q ~	[q ~�q ~�q ~bxq ~�sq ~`w    ?@     q ~ �q ~�q ~�q ~�q ~2q ~rq ~	=q ~1q ~�q ~q ~�q ~;q ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�q ~�q ~ q ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�xxsq ~ J?@     w       q ~5sq ~`w   ?@     q ~0q ~�xq ~�sq ~`w   @?@     *q ~Aq ~Vq ~�q ~q ~/q ~�q ~2q ~Nq ~�q ~
]q ~xq ~	�q ~$q ~�q ~^q ~�q ~�q ~q ~
q ~Sq ~q ~Gq ~	�q ~�q ~bq ~�q ~xq ~uq ~�q ~0q ~{q ~	�q ~�q ~�q ~�q ~	�q ~lq ~�q ~Jq ~{q ~Xq ~�xq ~
�sq ~`w   ?@     q ~
�xq ~�sq ~`w    ?@     q ~[q ~tq ~�q ~�q ~nq ~*q ~�q ~�q ~�q ~
iq ~�q ~q ~
q ~�q ~7q ~Dq ~q ~$q ~,q ~Vxq ~�sq ~`w   ?@     q ~�q ~jq ~�q ~�xq ~�sq ~`w   ?@     q ~�xq ~[sq ~`w   ?@     q ~Vxq ~vsq ~`w   ?@     q ~qxq ~�sq ~`w   ?@     q ~�q ~�q ~�xq ~tsq ~`w   ?@     q ~oxq ~�sq ~`w   ?@     q ~�xq ~csq ~`w   ?@     q ~�q ~�q ~uq ~�q ~^xq ~�sq ~`w   ?@     q ~�q ~�q ~�q ~	mq ~�q ~q ~
2q ~�xq ~�sq ~`w   ?@     
q ~
�q ~ q ~�q ~�q ~-q ~
�q ~q ~�q ~q ~�xq ~�sq ~`w   ?@     q ~�xq ~�sq ~`w   ?@     q ~�xq ~Csq ~`w   ?@     q ~�q ~>xq ~�sq ~`w   ?@     q ~<q ~�q ~�q ~�xq ~�sq ~`w   ?@     q ~�q ~	xq ~hsq ~`w   ?@     q ~cxxsr 9edu.cornell.cs.nlp.spf.base.hashvector.FastTreeHashVector;��tQ57� L valuest 0Lit/unimi/dsi/fastutil/objects/Object2DoubleMap;xpsr 5it.unimi.dsi.fastutil.objects.Object2DoubleAVLTreeMap�7y�J| I countL storedComparatort Ljava/util/Comparator;xr <it.unimi.dsi.fastutil.objects.AbstractObject2DoubleSortedMap�c����  xr 6it.unimi.dsi.fastutil.objects.AbstractObject2DoubleMap�o��K<z  xr ;it.unimi.dsi.fastutil.objects.AbstractObject2DoubleFunction�o��K<z D defRetValuexp          �psq ~mWD�t DYNSKIPppppw��      sq ~mW�"�q ~ t LEXt 0t 0pw        sq ~mW���q ~ q ~t 0t 22pw@$      sq ~mW��aq ~ q ~t 0t 39pw@$      sq ~mW�#�q ~ q ~t 0t 7pw        sq ~mW�&�q ~ q ~t 1t 1pw        sq ~mW���q ~ q ~t 1t 37pw@$      sq ~mW��
q ~ q ~t 1t 42pw        sq ~mW�!q ~ q ~t 10t 11pw        sq ~mW�iDq ~ q ~t 10t 2pw@@�鹙�sq ~mZw,�q ~ q ~t 100t 15pw@$      sq ~mZw0Hq ~ q ~t 100t 22pw        sq ~mZ�v9q ~ q ~t 101t 110pw@$      sq ~mZwC�q ~ q ~t 101t 66pw        sq ~mZwGJq ~ q ~t 101t 76pw@$      sq ~mZ�y�q ~ q ~t 102t 110pw@$      sq ~mZwGJq ~ q ~t 102t 66pw        sq ~mZwKq ~ q ~t 102t 76pw@$      sq ~mZwG+q ~ q ~t 103t 55pw@$      sq ~mZwRnq ~ q ~t 103t 85pw        sq ~mZwNq ~ q ~t 104t 60pw@$      sq ~mZwQ�q ~ q ~t 105t 60pw@$      sq ~mZ���q ~ q ~t 106t 110pw@$      sq ~mZwY�q ~ q ~t 106t 72pw        sq ~mZwZq ~ q ~t 106t 76pw@$      sq ~mZwa�q ~ q ~t 107t 86pw@5oz�G�sq ~mZ���q ~ q ~t 108t 110pw@$      sq ~mZw]�q ~ q ~t 108t 66pw        sq ~mZwa�q ~ q ~t 108t 76pw@$      sq ~mZwi2q ~ q ~t 109t 87pw@$      sq ~mZwl�q ~ q ~t 109t 94pw@$      sq ~mW�%q ~ q ~t 11t 13pw@$      sq ~mW�;>q ~ q ~t 11t 70pw@$      sq ~mW�m�q ~ q ~t 11t 9pw        sq ~mW�B�q ~ q ~t 11t 90pw@$      sq ~mZw��q ~ q ~t 110t 88pw        sq ~mZw��q ~ q ~t 110t 98pw@$      sq ~mZ��q ~ q ~t 111t 110pw@$      sq ~mZw��q ~ q ~t 111t 66pw        sq ~mZw��q ~ q ~t 111t 76pw@$      sq ~mZwq ~ q ~t 112t 81pw@5oz�G�sq ~mZwÈq ~ q ~t 112t 89pw        sq ~mZw��q ~ q ~t 112t 96pw@5oz�G�sq ~mZw��q ~ q ~t 113t 17pw        sq ~mZw��q ~ q ~t 113t 43pw@$      sq ~mZw�q ~ q ~t 113t 63pw@$      sq ~mZw�qq ~ q ~t 114t 60pw@$      sq ~mZ���q ~ q ~t 115t 110pw@$      sq ~mZw��q ~ q ~t 115t 66pw        sq ~mZw�1q ~ q ~t 115t 72pw@$      sq ~mZ���q ~ q ~t 116t 100pw@$      sq ~mZw��q ~ q ~t 116t 67pw        sq ~mZ�q ~ q ~t 117t 110pw@$      sq ~mZw�nq ~ q ~t 117t 66pw        sq ~mZw�/q ~ q ~t 117t 76pw@$      sq ~mZ��q ~ q ~t 118t 110pw@$      sq ~mZw�/q ~ q ~t 118t 66pw        sq ~mZw��q ~ q ~t 118t 76pw@$      sq ~mZw�q ~ q ~t 119t 83pw@5oz�G�sq ~mZw�q ~ q ~t 119t 92pw@5oz�G�sq ~mW�(�q ~ q ~t 12t 12pw        sq ~mW�4�q ~ q ~t 12t 48pw@$      sq ~mZx/mq ~ q ~t 120t 81pw@$      sq ~mZx3lq ~ q ~t 120t 93pw        sq ~mZx3�q ~ q ~t 120t 96pw@$      sq ~mZx3.q ~ q ~t 121t 81pw@$      sq ~mZx4&q ~ q ~t 121t 89pw        sq ~mZx7�q ~ q ~t 121t 96pw@$      sq ~mZx;,q ~ q ~t 122t 95pw        sq ~mZx;�q ~ q ~t 122t 98pw@$      sq ~mZx3q ~ q ~t 123t 60pw@$      sq ~mZx6�q ~ q ~t 124t 60pw@$      sq ~mZx/Nq ~ q ~t 125t 30pw@$      sq ~mZx0Fq ~ q ~t 125t 38pw        sq ~mZx>Rq ~ q ~t 126t 60pw@$      sq ~mZx7-q ~ q ~t 127t 33pw@$      sq ~mZx7�q ~ q ~t 127t 38pw        sq ~mZxNNq ~ q ~t 128t 88pw@$      sq ~mZxQ�q ~ q ~t 128t 95pw        sq ~mZxRq ~ q ~t 128t 98pw@$      sq ~mZxQ�q ~ q ~t 129t 87pw@5oz�G�sq ~mZxU5q ~ q ~t 129t 93pw        sq ~mZxUTq ~ q ~t 129t 94pw@5oz�G�sq ~mZxU�q ~ q ~t 129t 96pw        sq ~mW�,�q ~ q ~t 13t 13pw        sq ~mW�?\q ~ q ~t 13t 63pw@5oz�G�sq ~mW�@q ~ q ~t 13t 69pw        sq ~mZ�ϕq ~ q ~t 130t 110pw@$      sq ~mZx��q ~ q ~t 130t 66pw        sq ~mZx��q ~ q ~t 130t 76pw@$      sq ~mZ��Vq ~ q ~t 131t 110pw@$      sq ~mZx�gq ~ q ~t 131t 76pw@$      sq ~mZ��q ~ q ~t 132t 110pw@$      sq ~mZx��q ~ q ~t 132t 72pw        sq ~mZx�(q ~ q ~t 132t 76pw@$      sq ~mZx�nq ~ q ~t 133t 60pw@5oz�G�sq ~mZx�/q ~ q ~t 134t 60pw@$      sq ~mZx��q ~ q ~t 135t 83pw@$      sq ~mZx�qq ~ q ~t 135t 92pw@$      sq ~mZ��q ~ q ~t 136t 110pw@$      sq ~mZx��q ~ q ~t 136t 72pw        sq ~mZx�,q ~ q ~t 136t 76pw@$      sq ~mZ���q ~ q ~t 137t 110pw@5oz�G�sq ~mZx�qq ~ q ~t 137t 72pw@5oz�G�sq ~mZx�3q ~ q ~t 138t 60pw@$      sq ~mZx��q ~ q ~t 139t 60pw@$      sq ~mW�0wq ~ q ~t 14t 14pw        sq ~mW�3�q ~ q ~t 14t 20pw@$      sq ~mZ�C�q ~ q ~t 140t 110pw@$      sq ~mZyDq ~ q ~t 140t 66pw        sq ~mZyq ~ q ~t 140t 76pw@$      sq ~mZy gq ~ q ~t 141t 97pw@@�鹙�sq ~mZ�Kvq ~ q ~t 142t 110pw@$      sq ~mZyq ~ q ~t 142t 72pw        sq ~mZy�q ~ q ~t 142t 76pw@$      sq ~mZ�O7q ~ q ~t 143t 110pw@5oz�G�sq ~mZy�q ~ q ~t 143t 66pw        sq ~mZy Hq ~ q ~t 143t 76pw@5oz�G�sq ~mZ�R�q ~ q ~t 144t 110pw@$      sq ~mZy Hq ~ q ~t 144t 66pw        sq ~mZy#�q ~ q ~t 144t 72pw@$      sq ~mZy/�q ~ q ~t 145t 99pw@$      sq ~mZ�Zzq ~ q ~t 146t 110pw@5oz�G�sq ~mZy+q ~ q ~t 146t 72pw@5oz�G�sq ~mZy+�q ~ q ~t 146t 76pw        sq ~mZ�^;q ~ q ~t 147t 110pw@$      sq ~mZy+�q ~ q ~t 147t 66pw        sq ~mZy/Lq ~ q ~t 147t 76pw@$      sq ~mZy:pq ~ q ~t 148t 95pw@$      sq ~mZy:�q ~ q ~t 148t 98pw@$      sq ~mZy2Sq ~ q ~t 149t 60pw@$      sq ~mW�{�q ~ q ~t 15t 0pw        sq ~mW�7�q ~ q ~t 15t 22pw        sq ~mW�>�q ~ q ~t 15t 40pw@$      sq ~mZy��q ~ q ~t 150t 60pw@$      sq ~mZy�dq ~ q ~t 151t 66pw        sq ~mZy�%q ~ q ~t 151t 76pw@@�鹙�sq ~mZ���q ~ q ~t 152t 110pw@$      sq ~mZy�jq ~ q ~t 152t 72pw@$      sq ~mZy��q ~ q ~t 152t 76pw        sq ~mZy��q ~ q ~t 153t 66pw@@�鹙�sq ~mZy��q ~ q ~t 153t 76pw        sq ~mZ��Wq ~ q ~t 154t 110pw@$      sq ~mZy�hq ~ q ~t 154t 76pw@$      sq ~mZy��q ~ q ~t 155t 60pw@$      sq ~mZy�Hq ~ q ~t 156t 67pw        sq ~mZy��q ~ q ~t 156t 73pw@$      sq ~mZy��q ~ q ~t 156t 74pw@$      sq ~mZ���q ~ q ~t 157t 101pw@5oz�G�sq ~mZ���q ~ q ~t 157t 109pw@5oz�G�sq ~mZ��[q ~ q ~t 158t 110pw@F�U�i�sq ~mZy��q ~ q ~t 158t 72pw@F�U�i�sq ~mZy�lq ~ q ~t 158t 76pw        sq ~mZ��q ~ q ~t 159t 110pw@$      sq ~mZy��q ~ q ~t 159t 72pw        sq ~mZy�-q ~ q ~t 159t 76pw@$      sq ~mW�8q ~ q ~t 16t 15pw        sq ~mWĀ�q ~ q ~t 16t 8pw@$      sq ~mZ�,�q ~ q ~t 160t 110pw@$      sq ~mZy��q ~ q ~t 160t 76pw@$      sq ~mZy�	q ~ q ~t 161t 60pw@$      sq ~mZz �q ~ q ~t 162t 60pw@$      sq ~mZz�q ~ q ~t 163t 60pw@$      sq ~mZzLq ~ q ~t 164t 60pw@5oz�G�sq ~mZ�;�q ~ q ~t 165t 102pw@$      sq ~mZ�<Qq ~ q ~t 165t 105pw@$      sq ~mZ�?�q ~ q ~t 166t 103pw@5oz�G�sq ~mZ�F�q ~ q ~t 167t 110pw@$      sq ~mZz�q ~ q ~t 167t 72pw@$      sq ~mZzPq ~ q ~t 168t 60pw@$      sq ~mZzq ~ q ~t 169t 60pw@$      sq ~mW�;�q ~ q ~t 17t 16pw        sq ~mW�?�q ~ q ~t 17t 28pw@$      sq ~mW�Jaq ~ q ~t 17t 51pw@$      sq ~mZ��q ~ q ~t 170t 110pw@$      sq ~mZzq�q ~ q ~t 170t 72pw        sq ~mZzr"q ~ q ~t 170t 76pw@$      sq ~mZzqhq ~ q ~t 171t 60pw@5oz�G�sq ~mZz}q ~ q ~t 172t 83pw@$      sq ~mZz��q ~ q ~t 172t 92pw@$      sq ~mZ��Tq ~ q ~t 173t 110pw@$      sq ~mZzy�q ~ q ~t 173t 66pw        sq ~mZz}eq ~ q ~t 173t 76pw@$      sq ~mZz|�q ~ q ~t 174t 60pw@@�鹙�sq ~mZ���q ~ q ~t 175t 110pw@$      sq ~mZz�kq ~ q ~t 175t 72pw@$      sq ~mZ��Rq ~ q ~t 176t 104pw@5oz�G�sq ~mZz��q ~ q ~t 177t 60pw@$      sq ~mZz��q ~ q ~t 178t 60pw@$      sq ~mZz�pq ~ q ~t 179t 60pw@$      sq ~mW�?q ~ q ~t 18t 11pw@$      sq ~mW�?=q ~ q ~t 18t 12pw        sq ~mW�C�q ~ q ~t 18t 28pw        sq ~mZz��q ~ q ~t 180t 83pw@5oz�G�sq ~mZz�q ~ q ~t 180t 92pw@5oz�G�sq ~mZz��q ~ q ~t 181t 60pw@$      sq ~mZz�q ~ q ~t 182t 60pw@5oz�G�sq ~mZ� �q ~ q ~t 183t 110pw@$      sq ~mZz�Hq ~ q ~t 183t 72pw        sq ~mZz��q ~ q ~t 183t 76pw@$      sq ~mZz�
q ~ q ~t 184t 60pw@$      sq ~mZ�%.q ~ q ~t 185t 106pw@@�鹙�sq ~mZ�)q ~ q ~t 186t 107pw@5oz�G�sq ~mZz�Mq ~ q ~t 187t 60pw@$      sq ~mZ{ q ~ q ~t 188t 60pw@F�U�i�sq ~mZ{�q ~ q ~t 189t 60pw@$      sq ~mW�C�q ~ q ~t 19t 17pw        sq ~mW�F�q ~ q ~t 19t 21pw        sq ~mW�Vq ~ q ~t 19t 64pw@$      sq ~mW�V�q ~ q ~t 19t 69pw@$      sq ~mWċ�q ~ q ~t 19t 9pw@$      sq ~mZ��q ~ q ~t 190t 108pw@@�鹙�sq ~mZ{Z&q ~ q ~t 191t 60pw@$      sq ~mZ{]�q ~ q ~t 192t 60pw@$      sq ~mZ{a�q ~ q ~t 193t 60pw@5oz�G�sq ~mZ{eiq ~ q ~t 194t 60pw@$      sq ~mZ{i*q ~ q ~t 195t 60pw@$      sq ~mZ{l�q ~ q ~t 196t 60pw@$      sq ~mW�*xq ~ q ~t 2t 1pw@$      sq ~mW�*�q ~ q ~t 2t 2pw        sq ~mW��q ~ q ~t 2t 24pw        sq ~mWŖNq ~ q ~t 20t 18pw        sq ~mWŝ5q ~ q ~t 20t 33pw@$      sq ~mWŠ�q ~ q ~t 20t 43pw        sq ~mWšq ~ q ~t 20t 44pw        sq ~mWŤ�q ~ q ~t 20t 52pw        sq ~mWū�q ~ q ~t 20t 70pw        sq ~mWŬ�q ~ q ~t 20t 77pw@$      sq ~mWų^q ~ q ~t 20t 90pw        sq ~mWř�q ~ q ~t 21t 14pw@$      sq ~mWř�q ~ q ~t 21t 15pw        sq ~mWŝ�q ~ q ~t 22t 19pw        sq ~mWŬXq ~ q ~t 22t 54pw@$      sq ~mWŤZq ~ q ~t 23t 20pw        sq ~mWū�q ~ q ~t 23t 41pw@$      sq ~mW��iq ~ q ~t 24t 0pw@$      sq ~mWŨxq ~ q ~t 24t 23pw        sq ~mWŴVq ~ q ~t 24t 58pw        sq ~mWŨ�q ~ q ~t 25t 17pw        sq ~mWũq ~ q ~t 25t 18pw@$      sq ~mWů�q ~ q ~t 25t 30pw@$      sq ~mWů�q ~ q ~t 25t 33pw@$      sq ~mWŷq ~ q ~t 25t 50pw@$      sq ~mW���q ~ q ~t 25t 6pw@$      sq ~mWſzq ~ q ~t 25t 77pw@$      sq ~mWŬ�q ~ q ~t 26t 19pw        sq ~mWŻ�q ~ q ~t 26t 58pw@$      sq ~mWų�q ~ q ~t 27t 24pw@$      sq ~mWų�q ~ q ~t 27t 25pw        sq ~mWŻ{q ~ q ~t 27t 45pw        sq ~mW���q ~ q ~t 28t 100pw        sq ~mWŷ�q ~ q ~t 28t 26pw@@�鹙�sq ~mWŻ�q ~ q ~t 29t 27pw@$      sq ~mW�ƀq ~ q ~t 29t 53pw@$      sq ~mW���q ~ q ~t 29t 56pw@$      sq ~mW��@q ~ q ~t 29t 75pw@$      sq ~mW�.wq ~ q ~t 3t 3pw        sq ~mW��Gq ~ q ~t 3t 36pw@$      sq ~mW�	�q ~ q ~t 30t 10pw        sq ~mW��q ~ q ~t 30t 35pw@5oz�G�sq ~mW�R@q ~ q ~t 30t 4pw@5oz�G�sq ~mW�Vq ~ q ~t 31t 21pw        sq ~mW� �q ~ q ~t 31t 63pw        sq ~mW� �q ~ q ~t 31t 64pw        sq ~mW�!Rq ~ q ~t 31t 69pw@5oz�G�sq ~mW�Z]q ~ q ~t 32t 9pw        sq ~mW�/?q ~ q ~t 32t 90pw@$      sq ~mW��q ~ q ~t 33t 31pw@$      sq ~mW�]�q ~ q ~t 33t 5pw        sq ~mW��q ~ q ~t 34t 29pw        sq ~mW�%q ~ q ~t 34t 49pw        sq ~mW�(9q ~ q ~t 34t 54pw        sq ~mW�a�q ~ q ~t 34t 7pw@$      sq ~mW�#�q ~ q ~t 35t 30pw        sq ~mW�+�q ~ q ~t 35t 52pw@$      sq ~mW�'�q ~ q ~t 36t 30pw        sq ~mW�+�q ~ q ~t 36t 43pw@$      sq ~mW�/?q ~ q ~t 36t 50pw        sq ~mW�3]q ~ q ~t 36t 63pw@$      sq ~mW�>Cq ~ q ~t 36t 90pw@$      sq ~mW�+�q ~ q ~t 37t 31pw        sq ~mW�,Wq ~ q ~t 37t 37pw        sq ~mW�6�q ~ q ~t 37t 61pw@F�U�i�sq ~mW�,Wq ~ q ~t 38t 27pw@$      sq ~mW�/}q ~ q ~t 38t 32pw        sq ~mW�,Wq ~ q ~t 39t 17pw@$      sq ~mW�,vq ~ q ~t 39t 18pw@$      sq ~mW�3 q ~ q ~t 39t 30pw@$      sq ~mW�3]q ~ q ~t 39t 33pw        sq ~mW�2Wq ~ q ~t 4t 4pw        sq ~mW���q ~ q ~t 4t 51pw        sq ~mW��,q ~ q ~t 4t 65pw@$      sq ~mWƆq ~ q ~t 40t 34pw@$      sq ~mW��"q ~ q ~t 41t 2pw@$      sq ~mWƉ�q ~ q ~t 41t 35pw        sq ~mWƍ�q ~ q ~t 42t 36pw        sq ~mWƑ�q ~ q ~t 42t 49pw@$      sq ~mWƘ�q ~ q ~t 42t 65pw        sq ~mWƑ�q ~ q ~t 43t 38pw        sq ~mW��}q ~ q ~t 43t 9pw@5oz�G�sq ~mWƍq ~ q ~t 44t 10pw@$      sq ~mWƕ�q ~ q ~t 44t 39pw        sq ~mWƑq ~ q ~t 45t 12pw@$      sq ~mWƜq ~ q ~t 45t 40pw        sq ~mWƟ�q ~ q ~t 46t 41pw        sq ~mWƠxq ~ q ~t 46t 45pw@$      sq ~mWƘ�q ~ q ~t 47t 15pw@5oz�G�sq ~mWƜq ~ q ~t 47t 20pw        sq ~mWƠ:q ~ q ~t 48t 23pw@$      sq ~mWƤq ~ q ~t 48t 34pw        sq ~mWƫ^q ~ q ~t 49t 42pw        sq ~mWƲ�q ~ q ~t 49t 61pw@$      sq ~mW��Fq ~ q ~t 5t 28pw@$      sq ~mW�67q ~ q ~t 5t 5pw        sq ~mW��3q ~ q ~t 50t 32pw@5oz�G�sq ~mW��q ~ q ~t 50t 82pw@5oz�G�sq ~mW�Pq ~ q ~t 51t 47pw        sq ~mW��q ~ q ~t 51t 78pw@$      sq ~mW���q ~ q ~t 52t 29pw@$      sq ~mW��q ~ q ~t 52t 34pw        sq ~mW�	7q ~ q ~t 53t 42pw@$      sq ~mW�	�q ~ q ~t 53t 48pw        sq ~mW��q ~ q ~t 53t 62pw        sq ~mW��q ~ q ~t 54t 12pw        sq ~mW�q ~ q ~t 54t 15pw@5oz�G�sq ~mW�	q ~ q ~t 55t 21pw        sq ~mW�q ~ q ~t 55t 69pw@5oz�G�sq ~mW��q ~ q ~t 56t 27pw@$      sq ~mW��q ~ q ~t 56t 32pw@$      sq ~mW�Zq ~ q ~t 56t 53pw        sq ~mW� q ~ q ~t 56t 75pw        sq ~mW�#~q ~ q ~t 56t 82pw@$      sq ~mW��q ~ q ~t 57t 22pw@$      sq ~mW�Udq ~ q ~t 57t 5pw        sq ~mW� q ~ q ~t 58t 55pw        sq ~mW�+]q ~ q ~t 58t 85pw@$      sq ~mW�.�q ~ q ~t 58t 91pw@$      sq ~mW��q ~ q ~t 59t 27pw@$      sq ~mW��q ~ q ~t 59t 32pw@$      sq ~mW�#�q ~ q ~t 59t 56pw        sq ~mW�.�q ~ q ~t 59t 82pw@$      sq ~mW�.�q ~ q ~t 59t 84pw        sq ~mW�:q ~ q ~t 6t 6pw        sq ~mW�Vq ~ q ~t 6t 90pw@5oz�G�sq ~mW�klq ~ q ~t 60t 27pw@$      sq ~mW�v�q ~ q ~t 60t 59pw        sq ~mW�}Xq ~ q ~t 61t 60pw@$      sq ~mW�y�q ~ q ~t 62t 41pw        sq ~mWǁWq ~ q ~t 62t 62pw@5oz�G�sq ~mW�~q ~ q ~t 63t 46pw@$      sq ~mWǄ�q ~ q ~t 63t 61pw        sq ~mW�zpq ~ q ~t 64t 27pw        sq ~mW�}�q ~ q ~t 64t 32pw@$      sq ~mWǐ[q ~ q ~t 64t 82pw@$      sq ~mWǌ\q ~ q ~t 65t 60pw@$      sq ~mWǁ�q ~ q ~t 66t 26pw        sq ~mWǔ;q ~ q ~t 66t 73pw@$      sq ~mW��Hq ~ q ~t 67t 110pw@$      sq ~mWǔ�q ~ q ~t 67t 66pw        sq ~mWǘYq ~ q ~t 67t 76pw@$      sq ~mWǘxq ~ q ~t 68t 67pw@5oz�G�sq ~mWǌ{q ~ q ~t 69t 21pw@$      sq ~mWǜXq ~ q ~t 69t 68pw        sq ~mW�={q ~ q ~t 7t 3pw@$      sq ~mW�>q ~ q ~t 7t 8pw        sq ~mW��Tq ~ q ~t 70t 51pw        sq ~mW��q ~ q ~t 70t 57pw@$      sq ~mW���q ~ q ~t 71t 34pw        sq ~mW�'�q ~ q ~t 71t 5pw@$      sq ~mW��mq ~ q ~t 72t 16pw@$      sq ~mW��Lq ~ q ~t 72t 39pw        sq ~mW��q ~ q ~t 73t 19pw@5oz�G�sq ~mW���q ~ q ~t 73t 41pw        sq ~mW� �q ~ q ~t 74t 71pw        sq ~mW�|q ~ q ~t 74t 80pw@$      sq ~mW��qq ~ q ~t 75t 26pw        sq ~mW��q ~ q ~t 75t 73pw@$      sq ~mW��1q ~ q ~t 76t 38pw        sq ~mW�:�q ~ q ~t 76t 6pw@$      sq ~mW���q ~ q ~t 77t 13pw        sq ~mW��q ~ q ~t 77t 77pw        sq ~mW�>�q ~ q ~t 77t 9pw@5oz�G�sq ~mW��Pq ~ q ~t 78t 19pw        sq ~mW���q ~ q ~t 78t 25pw@$      sq ~mW��q ~ q ~t 79t 27pw@$      sq ~mW�[q ~ q ~t 79t 53pw        sq ~mW�Jq ~ q ~t 8t 38pw@$      sq ~mW��q ~ q ~t 8t 44pw@$      sq ~mW�A�q ~ q ~t 8t 6pw@$      sq ~mW��q ~ q ~t 8t 68pw@$      sq ~mW�A�q ~ q ~t 8t 9pw        sq ~mWޕ�q ~ q ~t 80t 110pw@5oz�G�sq ~mW�fTq ~ q ~t 80t 72pw@5oz�G�sq ~mW�W�q ~ q ~t 81t 27pw@$      sq ~mW�_mq ~ q ~t 81t 47pw@$      sq ~mW�cq ~ q ~t 81t 56pw@$      sq ~mW�jrq ~ q ~t 81t 75pw@$      sq ~mW�nq ~ q ~t 81t 84pw@$      sq ~mWޝAq ~ q ~t 82t 110pw@$      sq ~mW�m�q ~ q ~t 82t 72pw        sq ~mW�nRq ~ q ~t 82t 76pw@$      sq ~mW�jrq ~ q ~t 83t 55pw        sq ~mW�u�q ~ q ~t 83t 86pw@$      sq ~mW�_�q ~ q ~t 84t 18pw@$      sq ~mW�fq ~ q ~t 84t 30pw@$      sq ~mW�q�q ~ q ~t 84t 64pw        sq ~mW�y8q ~ q ~t 85t 73pw@$      sq ~mW�yWq ~ q ~t 85t 74pw@$      sq ~mWެEq ~ q ~t 86t 110pw@$      sq ~mW�}Vq ~ q ~t 86t 76pw@$      sq ~mW�q�q ~ q ~t 87t 32pw@5oz�G�sq ~mWȁUq ~ q ~t 87t 78pw        sq ~mWȄ\q ~ q ~t 87t 82pw@5oz�G�sq ~mWȀ]q ~ q ~t 88t 60pw@$      sq ~mWȈ�q ~ q ~t 89t 79pw@@�鹙�sq ~mW���q ~ q ~t 9t 10pw        sq ~mW�2q ~ q ~t 9t 31pw@5oz�G�sq ~mW��q ~ q ~t 9t 46pw        sq ~mW�nq ~ q ~t 9t 57pw        sq ~mW�ȉq ~ q ~t 90t 27pw@$      sq ~mW�ӭq ~ q ~t 90t 56pw        sq ~mW��
q ~ q ~t 90t 59pw@$      sq ~mW���q ~ q ~t 91t 80pw        sq ~mW��q ~ q ~t 91t 89pw@@�鹙�sq ~mW��4q ~ q ~t 91t 94pw        sq ~mW��q ~ q ~t 92t 110pw@$      sq ~mW��5q ~ q ~t 92t 72pw        sq ~mW��q ~ q ~t 92t 76pw@$      sq ~mW�aq ~ q ~t 93t 110pw@5oz�G�sq ~mW��q ~ q ~t 93t 66pw        sq ~mW���q ~ q ~t 93t 72pw@5oz�G�sq ~mW��q ~ q ~t 94t 71pw@5oz�G�sq ~mW��Yq ~ q ~t 94t 81pw        sq ~mW��Xq ~ q ~t 94t 93pw@5oz�G�sq ~mW��Nq ~ q ~t 95t 27pw@$      sq ~mW���q ~ q ~t 95t 59pw@$      sq ~mW���q ~ q ~t 95t 75pw        sq ~mW� �q ~ q ~t 96t 110pw@$      sq ~mW��9q ~ q ~t 96t 72pw        sq ~mW��q ~ q ~t 96t 76pw@$      sq ~mW���q ~ q ~t 97t 83pw@$      sq ~mW��|q ~ q ~t 97t 92pw@$      sq ~mW�(&q ~ q ~t 98t 110pw@$      sq ~mW���q ~ q ~t 98t 72pw        sq ~mW��7q ~ q ~t 98t 76pw@$      sq ~mW�+�q ~ q ~t 99t 110pw@$      sq ~mW��7q ~ q ~t 99t 66pw        sq ~mW��|q ~ q ~t 99t 72pw@$      q ~rw?�      sq ~me��q ~ t TMPt 0ppw        sq ~me���q ~ q ~?t 1ppw        sq ~me�A>q ~ q ~?t 10ppw        sq ~mh�L�q ~ q ~?t 100ppw        sq ~mh�PQq ~ q ~?t 101ppw        sq ~mh�Tq ~ q ~?t 102ppw        sq ~mh�W�q ~ q ~?t 103ppw        sq ~mh�[�q ~ q ~?t 104ppw        sq ~mh�_Uq ~ q ~?t 105ppw        sq ~mh�cq ~ q ~?t 106ppw        sq ~mh�f�q ~ q ~?t 107ppw        sq ~mh�j�q ~ q ~?t 108ppw        sq ~mh�nYq ~ q ~?t 109ppw        sq ~me�D�q ~ q ~?t 11ppw        sq ~mh���q ~ q ~?t 110ppw        sq ~me�H�q ~ q ~?t 12ppw        sq ~me�L�q ~ q ~?t 13ppw        sq ~me�PBq ~ q ~?t 14ppw        sq ~me�Tq ~ q ~?t 15ppw        sq ~me�W�q ~ q ~?t 16ppw        sq ~me�[�q ~ q ~?t 17ppw        sq ~me�_Fq ~ q ~?t 18ppw        sq ~me�cq ~ q ~?t 19ppw        sq ~me��q ~ q ~?t 2ppw        sq ~meص�q ~ q ~?t 20ppw        sq ~meع^q ~ q ~?t 21ppw        sq ~meؽq ~ q ~?t 22ppw        sq ~me���q ~ q ~?t 23ppw        sq ~me�ġq ~ q ~?t 24ppw        sq ~me��bq ~ q ~?t 25ppw        sq ~me��#q ~ q ~?t 26ppw        sq ~me���q ~ q ~?t 27ppw        sq ~me�ӥq ~ q ~?t 28ppw        sq ~me��fq ~ q ~?t 29ppw        sq ~me�Rq ~ q ~?t 3ppw        sq ~me�)�q ~ q ~?t 30ppw        sq ~me�-�q ~ q ~?t 31ppw        sq ~me�1~q ~ q ~?t 32ppw        sq ~me�5?q ~ q ~?t 33ppw        sq ~me�9 q ~ q ~?t 34ppw        sq ~me�<�q ~ q ~?t 35ppw        sq ~me�@�q ~ q ~?t 36ppw        sq ~me�DCq ~ q ~?t 37ppw        sq ~me�Hq ~ q ~?t 38ppw        sq ~me�K�q ~ q ~?t 39ppw        sq ~me�
q ~ q ~?t 4ppw        sq ~meٞ[q ~ q ~?t 40ppw        sq ~me٢q ~ q ~?t 41ppw        sq ~me٥�q ~ q ~?t 42ppw        sq ~me٩�q ~ q ~?t 43ppw        sq ~me٭_q ~ q ~?t 44ppw        sq ~meٱ q ~ q ~?t 45ppw        sq ~meٴ�q ~ q ~?t 46ppw        sq ~meٸ�q ~ q ~?t 47ppw        sq ~meټcq ~ q ~?t 48ppw        sq ~me��$q ~ q ~?t 49ppw        sq ~me��q ~ q ~?t 5ppw        sq ~me��q ~ q ~?t 50ppw        sq ~me�{q ~ q ~?t 51ppw        sq ~me�<q ~ q ~?t 52ppw        sq ~me��q ~ q ~?t 53ppw        sq ~me�!�q ~ q ~?t 54ppw        sq ~me�%q ~ q ~?t 55ppw        sq ~me�)@q ~ q ~?t 56ppw        sq ~me�-q ~ q ~?t 57ppw        sq ~me�0�q ~ q ~?t 58ppw        sq ~me�4�q ~ q ~?t 59ppw        sq ~me��q ~ q ~?t 6ppw        sq ~meڇq ~ q ~?t 60ppw        sq ~meڊ�q ~ q ~?t 61ppw        sq ~meڎ�q ~ q ~?t 62ppw        sq ~meڒ\q ~ q ~?t 63ppw        sq ~meږq ~ q ~?t 64ppw        sq ~meڙ�q ~ q ~?t 65ppw        sq ~meڝ�q ~ q ~?t 66ppw        sq ~meڡ`q ~ q ~?t 67ppw        sq ~meڥ!q ~ q ~?t 68ppw        sq ~meڨ�q ~ q ~?t 69ppw        sq ~me�Vq ~ q ~?t 7ppw        sq ~me��xq ~ q ~?t 70ppw        sq ~me��9q ~ q ~?t 71ppw        sq ~me��q ~ q ~?t 72ppw        sq ~me��q ~ q ~?t 73ppw        sq ~me�
|q ~ q ~?t 74ppw        sq ~me�=q ~ q ~?t 75ppw        sq ~me��q ~ q ~?t 76ppw        sq ~me��q ~ q ~?t 77ppw        sq ~me��q ~ q ~?t 78ppw        sq ~me�Aq ~ q ~?t 79ppw        sq ~me�q ~ q ~?t 8ppw        sq ~me�o�q ~ q ~?t 80ppw        sq ~me�s�q ~ q ~?t 81ppw        sq ~me�wYq ~ q ~?t 82ppw        sq ~me�{q ~ q ~?t 83ppw        sq ~me�~�q ~ q ~?t 84ppw        sq ~meۂ�q ~ q ~?t 85ppw        sq ~meۆ]q ~ q ~?t 86ppw        sq ~meۊq ~ q ~?t 87ppw        sq ~meۍ�q ~ q ~?t 88ppw        sq ~meۑ�q ~ q ~?t 89ppw        sq ~me��q ~ q ~?t 9ppw        sq ~me��6q ~ q ~?t 90ppw        sq ~me���q ~ q ~?t 91ppw        sq ~me��q ~ q ~?t 92ppw        sq ~me��yq ~ q ~?t 93ppw        sq ~me��:q ~ q ~?t 94ppw        sq ~me���q ~ q ~?t 95ppw        sq ~me���q ~ q ~?t 96ppw        sq ~me��}q ~ q ~?t 97ppw        sq ~me�>q ~ q ~?t 98ppw        sq ~me��q ~ q ~?t 99ppw        q ~nw?�      sq ~m{H�q ~ t XEMEt 0ppw@$      sq ~m{H��q ~ q ~t 1ppw@$      sq ~m{^�0q ~ q ~t 10ppw@$      sq ~m~��q ~ q ~t 100ppw@$      sq ~m~�Cq ~ q ~t 101ppw@$      sq ~m~q ~ q ~t 102ppw@$      sq ~m~�q ~ q ~t 103ppw@$      sq ~m~�q ~ q ~t 104ppw@$      sq ~m~Gq ~ q ~t 105ppw@$      sq ~m~q ~ q ~t 106ppw@$      sq ~m~�q ~ q ~t 107ppw@$      sq ~m~�q ~ q ~t 108ppw@$      sq ~m~Kq ~ q ~t 109ppw@$      sq ~m{^��q ~ q ~t 11ppw@$      sq ~m~m�q ~ q ~t 110ppw@$      sq ~m~q�q ~ q ~t 111ppw@$      sq ~m~ucq ~ q ~t 112ppw@$      sq ~m~y$q ~ q ~t 113ppw@$      sq ~m~|�q ~ q ~t 114ppw@$      sq ~m~��q ~ q ~t 115ppw@$      sq ~m~�gq ~ q ~t 116ppw@$      sq ~m~�(q ~ q ~t 117ppw@$      sq ~m~��q ~ q ~t 118ppw@$      sq ~m~��q ~ q ~t 119ppw@$      sq ~m{^��q ~ q ~t 12ppw@$      sq ~m~�@q ~ q ~t 120ppw@$      sq ~m~�q ~ q ~t 121ppw@$      sq ~m~��q ~ q ~t 122ppw@$      sq ~m~�q ~ q ~t 123ppw@$      sq ~m~�Dq ~ q ~t 124ppw@$      sq ~m~�q ~ q ~t 125ppw@$      sq ~m~��q ~ q ~t 126ppw@$      sq ~m~��q ~ q ~t 127ppw@$      sq ~m~ Hq ~ q ~t 128ppw@$      sq ~m~	q ~ q ~t 129ppw@$      sq ~m{^�sq ~ q ~t 13ppw@$      sq ~m~V�q ~ q ~t 130ppw@$      sq ~m~Z`q ~ q ~t 131ppw@$      sq ~m~^!q ~ q ~t 132ppw@$      sq ~m~a�q ~ q ~t 133ppw@$      sq ~m~e�q ~ q ~t 134ppw@$      sq ~m~idq ~ q ~t 135ppw@$      sq ~m~m%q ~ q ~t 136ppw@$      sq ~m~p�q ~ q ~t 137ppw@$      sq ~m~t�q ~ q ~t 138ppw@$      sq ~m~xhq ~ q ~t 139ppw@$      sq ~m{^�4q ~ q ~t 14ppw@$      sq ~m~��q ~ q ~t 140ppw@$      sq ~m~οq ~ q ~t 141ppw@$      sq ~m~Ҁq ~ q ~t 142ppw@$      sq ~m~�Aq ~ q ~t 143ppw@$      sq ~m~�q ~ q ~t 144ppw@$      sq ~m~��q ~ q ~t 145ppw@$      sq ~m~�q ~ q ~t 146ppw@$      sq ~m~�Eq ~ q ~t 147ppw@$      sq ~m~�q ~ q ~t 148ppw@$      sq ~m~��q ~ q ~t 149ppw@$      sq ~m{_ �q ~ q ~t 15ppw@$      sq ~m~?]q ~ q ~t 150ppw@$      sq ~m~Cq ~ q ~t 151ppw@$      sq ~m~F�q ~ q ~t 152ppw@$      sq ~m~J�q ~ q ~t 153ppw@$      sq ~m~Naq ~ q ~t 154ppw@$      sq ~m~R"q ~ q ~t 155ppw@$      sq ~m~U�q ~ q ~t 156ppw@$      sq ~m~Y�q ~ q ~t 157ppw@$      sq ~m~]eq ~ q ~t 158ppw@$      sq ~m~a&q ~ q ~t 159ppw@$      sq ~m{_�q ~ q ~t 16ppw@$      sq ~m~��q ~ q ~t 160ppw@$      sq ~m~�}q ~ q ~t 161ppw@$      sq ~m~�>q ~ q ~t 162ppw@$      sq ~m~��q ~ q ~t 163ppw@$      sq ~m~��q ~ q ~t 164ppw@$      sq ~m~Ɓq ~ q ~t 165ppw@$      sq ~m~�Bq ~ q ~t 166ppw@$      sq ~m~�q ~ q ~t 167ppw@$      sq ~m~��q ~ q ~t 168ppw@$      sq ~m~Յq ~ q ~t 169ppw@$      sq ~m{_wq ~ q ~t 17ppw@$      sq ~m~(q ~ q ~t 170ppw@$      sq ~m~+�q ~ q ~t 171ppw@$      sq ~m~/�q ~ q ~t 172ppw@$      sq ~m~3^q ~ q ~t 173ppw@$      sq ~m~7q ~ q ~t 174ppw@$      sq ~m~:�q ~ q ~t 175ppw@$      sq ~m~>�q ~ q ~t 176ppw@$      sq ~m~Bbq ~ q ~t 177ppw@$      sq ~m~F#q ~ q ~t 178ppw@$      sq ~m~I�q ~ q ~t 179ppw@$      sq ~m{_8q ~ q ~t 18ppw@$      sq ~m~�zq ~ q ~t 180ppw@$      sq ~m~�;q ~ q ~t 181ppw@$      sq ~m~��q ~ q ~t 182ppw@$      sq ~m~��q ~ q ~t 183ppw@$      sq ~m~�~q ~ q ~t 184ppw@$      sq ~m~�?q ~ q ~t 185ppw@$      sq ~m~� q ~ q ~t 186ppw@$      sq ~m~��q ~ q ~t 187ppw@$      sq ~m~��q ~ q ~t 188ppw@$      sq ~m~�Cq ~ q ~t 189ppw@$      sq ~m{_�q ~ q ~t 19ppw@$      sq ~m~�q ~ q ~t 190ppw@$      sq ~m~�q ~ q ~t 191ppw@$      sq ~m~[q ~ q ~t 192ppw@$      sq ~m~q ~ q ~t 193ppw@$      sq ~m~�q ~ q ~t 194ppw@$      sq ~m~#�q ~ q ~t 195ppw@$      sq ~m~'_q ~ q ~t 196ppw@$      sq ~m{H��q ~ q ~t 2ppw@$      sq ~m{_b�q ~ q ~t 20ppw@$      sq ~m{_fPq ~ q ~t 21ppw@$      sq ~m{_jq ~ q ~t 22ppw@$      sq ~m{_m�q ~ q ~t 23ppw@$      sq ~m{_q�q ~ q ~t 24ppw@$      sq ~m{_uTq ~ q ~t 25ppw@$      sq ~m{_yq ~ q ~t 26ppw@$      sq ~m{_|�q ~ q ~t 27ppw@$      sq ~m{_��q ~ q ~t 28ppw@$      sq ~m{_�Xq ~ q ~t 29ppw@$      sq ~m{H�Dq ~ q ~t 3ppw@$      sq ~m{_��q ~ q ~t 30ppw@$      sq ~m{_گq ~ q ~t 31ppw@$      sq ~m{_�pq ~ q ~t 32ppw@$      sq ~m{_�1q ~ q ~t 33ppw@$      sq ~m{_��q ~ q ~t 34ppw@$      sq ~m{_�q ~ q ~t 35ppw@$      sq ~m{_�tq ~ q ~t 36ppw@$      sq ~m{_�5q ~ q ~t 37ppw@$      sq ~m{_��q ~ q ~t 38ppw@$      sq ~m{_��q ~ q ~t 39ppw@$      sq ~m{H�q ~ q ~t 4ppw@$      sq ~m{`KMq ~ q ~t 40ppw@$      sq ~m{`Oq ~ q ~t 41ppw@$      sq ~m{`R�q ~ q ~t 42ppw@$      sq ~m{`V�q ~ q ~t 43ppw@$      sq ~m{`ZQq ~ q ~t 44ppw@$      sq ~m{`^q ~ q ~t 45ppw@$      sq ~m{`a�q ~ q ~t 46ppw@$      sq ~m{`e�q ~ q ~t 47ppw@$      sq ~m{`iUq ~ q ~t 48ppw@$      sq ~m{`mq ~ q ~t 49ppw@$      sq ~m{H��q ~ q ~t 5ppw@$      sq ~m{`��q ~ q ~t 50ppw@$      sq ~m{`�mq ~ q ~t 51ppw@$      sq ~m{`�.q ~ q ~t 52ppw@$      sq ~m{`��q ~ q ~t 53ppw@$      sq ~m{`ΰq ~ q ~t 54ppw@$      sq ~m{`�qq ~ q ~t 55ppw@$      sq ~m{`�2q ~ q ~t 56ppw@$      sq ~m{`��q ~ q ~t 57ppw@$      sq ~m{`ݴq ~ q ~t 58ppw@$      sq ~m{`�uq ~ q ~t 59ppw@$      sq ~m{H��q ~ q ~t 6ppw@$      sq ~m{a4q ~ q ~t 60ppw@$      sq ~m{a7�q ~ q ~t 61ppw@$      sq ~m{a;�q ~ q ~t 62ppw@$      sq ~m{a?Nq ~ q ~t 63ppw@$      sq ~m{aCq ~ q ~t 64ppw@$      sq ~m{aF�q ~ q ~t 65ppw@$      sq ~m{aJ�q ~ q ~t 66ppw@$      sq ~m{aNRq ~ q ~t 67ppw@$      sq ~m{aRq ~ q ~t 68ppw@$      sq ~m{aU�q ~ q ~t 69ppw@$      sq ~m{H�Hq ~ q ~t 7ppw@$      sq ~m{a�jq ~ q ~t 70ppw@$      sq ~m{a�+q ~ q ~t 71ppw@$      sq ~m{a��q ~ q ~t 72ppw@$      sq ~m{a��q ~ q ~t 73ppw@$      sq ~m{a�nq ~ q ~t 74ppw@$      sq ~m{a�/q ~ q ~t 75ppw@$      sq ~m{a��q ~ q ~t 76ppw@$      sq ~m{a±q ~ q ~t 77ppw@$      sq ~m{a�rq ~ q ~t 78ppw@$      sq ~m{a�3q ~ q ~t 79ppw@$      sq ~m{H�	q ~ q ~t 8ppw@$      sq ~m{b�q ~ q ~t 80ppw@$      sq ~m{b �q ~ q ~t 81ppw@$      sq ~m{b$Kq ~ q ~t 82ppw@$      sq ~m{b(q ~ q ~t 83ppw@$      sq ~m{b+�q ~ q ~t 84ppw@$      sq ~m{b/�q ~ q ~t 85ppw@$      sq ~m{b3Oq ~ q ~t 86ppw@$      sq ~m{b7q ~ q ~t 87ppw@$      sq ~m{b:�q ~ q ~t 88ppw@$      sq ~m{b>�q ~ q ~t 89ppw@$      sq ~m{H��q ~ q ~t 9ppw@$      sq ~m{b�(q ~ q ~t 90ppw@$      sq ~m{b��q ~ q ~t 91ppw@$      sq ~m{b��q ~ q ~t 92ppw@$      sq ~m{b�kq ~ q ~t 93ppw@$      sq ~m{b�,q ~ q ~t 94ppw@$      sq ~m{b��q ~ q ~t 95ppw@$      sq ~m{b��q ~ q ~t 96ppw@$      sq ~m{b�oq ~ q ~t 97ppw@$      sq ~m{b�0q ~ q ~t 98ppw@$      sq ~m{b��q ~ q ~t 99ppw@$      q ~pw?�      x