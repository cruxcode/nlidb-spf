�� sr -edu.cornell.cs.nlp.spf.parser.ccg.model.Model�5B��B�~ L featureSetst Ljava/util/List;L independentLexicalFeatureSetsq ~ L invalidFeaturest Ljava/util/Set;L lexicont -Ledu/cornell/cs/nlp/spf/ccg/lexicon/ILexicon;L thetat 4Ledu/cornell/cs/nlp/spf/base/hashvector/IHashVector;xpsr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.LinkedList)S]J`�"  xpw   sr Pedu.cornell.cs.nlp.spf.parser.ccg.factoredlex.features.FactoredLexicalFeatureSet�g�պ��� D 
entryScaleI lexemeNextIdD lexemeScaleI nonFactoredNextIdI templateNextIdD templateScaleL entryInitialScorert :Ledu/cornell/cs/nlp/utils/collections/ISerializableScorer;L 	lexemeIdst 5Lit/unimi/dsi/fastutil/objects/Object2IntOpenHashMap;L lexemeInitialScorerq ~ L nonFactoredIdsq ~ L templateIdsq ~ L templateInitialScorerq ~ xr Iedu.cornell.cs.nlp.spf.parser.ccg.model.lexical.AbstractLexicalFeatureSetZ���n3�� Z computeSyntaxAttributeFeaturesL 
featureTagt Ljava/lang/String;L ignoreFiltert Ljava/util/function/Predicate;xp t FACLEXsr !java.lang.invoke.SerializedLambdaoaД,)6� 
I implMethodKind[ capturedArgst [Ljava/lang/Object;L capturingClasst Ljava/lang/Class;L functionalInterfaceClassq ~ L functionalInterfaceMethodNameq ~ L "functionalInterfaceMethodSignatureq ~ L 	implClassq ~ L implMethodNameq ~ L implMethodSignatureq ~ L instantiatedMethodTypeq ~ xp   ur [Ljava.lang.Object;��X�s)l  xp    vr 0edu.cornell.cs.nlp.utils.function.PredicateUtils           xpt java/util/function/Predicatet testt (Ljava/lang/Object;)Zt 0edu/cornell/cs/nlp/utils/function/PredicateUtilst lambda$alwaysTrue$bcad8f2c$1q ~ q ~ ?�        
a?�             U?�������sr Eedu.cornell.cs.nlp.spf.parser.ccg.features.basic.scorer.UniformScorerQ�B���S D scorexp        sr 3it.unimi.dsi.fastutil.objects.Object2IntOpenHashMap         F fI sizexr 3it.unimi.dsi.fastutil.objects.AbstractObject2IntMap�o��K<z  xr 8it.unimi.dsi.fastutil.objects.AbstractObject2IntFunction�o��K<z I defRetValuexp    ?@    
asr 9edu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.Lexeme	I����� I hashCodeCacheL 
attributesq ~ L 	constantsq ~ L 
propertiest Ljava/util/Map;L 	signaturet GLedu/cornell/cs/nlp/spf/ccg/lexicon/factored/lambda/FactoringSignature;L tokenst ,Ledu/cornell/cs/nlp/spf/base/token/TokenSeq;xp`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sr 0edu.cornell.cs.nlp.spf.mr.lambda.LogicalConstant=Q��� L baseNameq ~ L nameq ~ xr %edu.cornell.cs.nlp.spf.mr.lambda.Term�(G^� L typet .Ledu/cornell/cs/nlp/spf/mr/language/type/Type;xr 2edu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression
n�tL�h  xpsr 0edu.cornell.cs.nlp.spf.mr.language.type.TermType��6��ǭ L parentt 2Ledu/cornell/cs/nlp/spf/mr/language/type/TermType;xr ,edu.cornell.cs.nlp.spf.mr.language.type.Typeg���� I hashCodeCacheL nameq ~ xp   st ssq ~ 5  �t losq ~ 5   et ept mainet maine:sxq ~ /q ~ .sr %java.util.Collections$UnmodifiableMap��t�B L mq ~ (xpsq ~ @sr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t origint fixed_domainxsr Eedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoringSignature�ڝ�U鞉 I hashCodeI numAttributesL typesq ~ xp  E    sq ~ sr java.util.ArrayListx����a� I sizexp   w   q ~ <xq ~ Ksr *edu.cornell.cs.nlp.spf.base.token.TokenSeq�py��An I hashCode[ tokenst [Ljava/lang/String;xpa��ur [Ljava.lang.String;��V��{G  xp   t thet statet ofq ~ >w  �sq ~ 'U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5   ct cq ~ :t dearborn_mit dearborn_mi:cxq ~ Xq ~ Wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ csq ~ LV0�uq ~ O   t dearbornt michiganw  �sq ~ '�<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5   mt mq ~ :t mount_evanst mount_evans:mxq ~ lq ~ ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ wsq ~ L��|uq ~ O   t mountt evansw  +sq ~ 'b=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5   rt rq ~ :t hudson_rivert hudson_river:rxq ~ �q ~ sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ LW��uq ~ O   q ~ Qt hudsont riverw  dsq ~ 'H��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sr 3edu.cornell.cs.nlp.spf.mr.language.type.ComplexType� �g��V L domainq ~ 2L rangeq ~ 2xq ~ 7=h��t <lo,<lo,t>>q ~ :sq ~ �l��Wt <lo,t>q ~ :sq ~ 5   tt tpt loct loc:<lo,<lo,t>>sq ~ 0q ~ 8t texast texas:sxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G��S    sq ~ sq ~ J   w   sq ~ �?z�t 	<e,<e,t>>q ~ <sq ~ �|-t <e,t>q ~ <q ~ �q ~ <xq ~ �sq ~ L�^�uq ~ O   q ~ �w   Hsq ~ '��|3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t bighorn_rivert bighorn_river:rxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L2�[�uq ~ O   t bighornq ~ �w   nsq ~ '�m�0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fort_smith_art fort_smith_ar:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L~�Suq ~ O   t fortt smitht arw  �sq ~ '�k(�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_bernardino_cat san_bernardino_ca:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L�Fuq ~ O   t sant 
bernardinot caw  sq ~ 'Unsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt el_cajon_cat el_cajon_ca:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L�w�uq ~ O   q ~ Qt cityt elt cajonw  osq ~ '0(�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_angelo_txt san_angelo_tx:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L&���uq ~ O   q ~ Qq ~ �q ~ �t angelow  usq ~ '�)M�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt salt_lake_city_utt salt_lake_city_ut:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L2�\Tuq ~ O   t saltt lakeq ~ �t utahw   �sq ~ 'Ҧ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 
californiat california:sxq ~ q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)sq ~ L:�M�uq ~ O   q ~ Qq ~ Rq ~ Sq ~"w  sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt portsmouth_vat portsmouth_va:cxq ~0q ~/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9sq ~ L�(6uq ~ O   t 
portsmoutht vaw   sq ~ '���<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t white_rivert white_river:rxq ~Bq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ksq ~ L��uq ~ O   q ~ Qt whitew   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt portland_ort portland_or:cxq ~Sq ~Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\sq ~ LC+MWuq ~ O   t portlandt orw  �sq ~ '�)��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt richmond_cat richmond_ca:cxq ~eq ~dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~nsq ~ L���duq ~ O   t richmondq ~"w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_york_cityt new_york_city:cxq ~vq ~usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��uq ~ O   t newt yorkt nyw  $sq ~ 'Ь��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5   nt nq ~ <t bellevuet 
bellevue:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lau��uq ~ O   q ~�w  |sq ~ '����sr java.util.Collections$EmptyListz��<���  xpsq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ ��|_t <s,t>q ~ 8q ~ �q ~ Rt state:<s,t>xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Et genlexxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ L��I�uq ~ O   t adjacentw  
Tsq ~ '���{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t little_rockt little_rock:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L_uq ~ O   t littlet rockw  Nsq ~ ')8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt providence_rit providence_ri:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L{(�uq ~ O   t 
providencet riw  �sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t mount_vernont mount_vernon:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�s�1uq ~ O   q ~ zt vernonw  	sq ~ 'n�$Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt des_moines_iat des_moines_ia:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�|�Cuq ~ O   t dest moinesw  �sq ~ 'N��Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
altoona_pat altoona_pa:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��̎uq ~ O   t altoonat pennsylvaniaw  �sq ~ '�ET�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
bristol_ctt bristol_ct:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L���uq ~ O   t bristolw   �sq ~ '�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t mobilet mobile:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"sq ~ L�J��uq ~ O   q ~w  Tsq ~ '�%�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t tennessee_rivert tennessee_river:rxq ~)q ~(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2sq ~ L�w%#uq ~ O   q ~ Qt 	tennesseew  sq ~ '�=�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt stockton_cat stockton_ca:cxq ~:q ~9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Csq ~ Lq��!uq ~ O   q ~ Qq ~ �t stocktonw  Msq ~ 'V�#rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t district_of_columbiat district_of_columbia:sxq ~Kq ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L�uq ~ O   q ~ Rq ~ St districtq ~ St columbiaw  Vsq ~ 'lg8}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~]q ~\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~csq ~ L%��duq ~ O   q ~ �q ~ �t arkansasw  	�sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	lawton_okt lawton_ok:cxq ~kq ~jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tsq ~ L��$�uq ~ O   t lawtonw  �sq ~ '�U�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t lawrencet 
lawrence:nxq ~|q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~~w  ]sq ~ '!�zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t marylandt 
maryland:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~�w  Ssq ~ '�#��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t normant norman:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��'uq ~ O   q ~�w  Esq ~ 'A�ݣsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t delawaret 
delaware:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�zuq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  %sq ~ '�tCzsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt youngstown_oht youngstown_oh:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   t 
youngstownw  }sq ~ '�R�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt las_vegas_nvt las_vegas_nv:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   t last vegasw  @sq ~ '��Xq ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ �t next_tot next_to:<lo,<lo,t>>xq ~�q ~�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ Luq ~ O   t bordersw  	�sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt daly_city_cat daly_city_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��suuq ~ O   t dalyq ~ �q ~"w  �sq ~ '�/Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bristol_township_pat bristol_township_pa:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LZw�Quq ~ O   q ~ Qq ~ �q ~t townshipw  �sq ~ '���6q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ �l��t <lo,i>q ~ :sq ~ 5   it iq ~ <t 
populationt population:<lo,i>xq ~q ~sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   sq ~ �|\t <e,e>q ~ <q ~ <xq ~sq ~ L  cuq ~ O   t inw  	�sq ~ '��4�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t los_angelest los_angeles:nxq ~#q ~"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,sq ~ L��R�uq ~ O   t lost angelesw   �sq ~ 'Z�X sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*xq ~5q ~4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;sq ~ LM�u�uq ~ O   q ~ Qq ~5q ~ �w  �sq ~ '�3vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t st_petersburgt st_petersburg:nxq ~Bq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ksq ~ L�uq ~ O   t stt 
petersburgw  sq ~ '<%�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt el_monte_cat el_monte_ca:cxq ~Tq ~Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]sq ~ L5��uq ~ O   q ~ �t montew  �sq ~ '��֠sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	tucson_azt tucson_az:cxq ~eq ~dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~nsq ~ L̑��uq ~ O   t tucsonw  Ssq ~ '&r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt charleston_wvt charleston_wv:cxq ~vq ~usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LF���uq ~ O   t 
charlestont wvw   �sq ~ 'qI��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt brockton_mat brockton_ma:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L"i�uq ~ O   q ~ Qq ~ �t brocktonw  �sq ~ ';E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���xuq ~ O   q ~ �q ~ �q ~ �w  �sq ~ '�?"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt ogden_utt 
ogden_ut:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Dq�uq ~ O   t ogdent utw  �sq ~ '��r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
alexandriat alexandria:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�8��uq ~ O   q ~�w  Tsq ~ '4=/�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cranston_rit cranston_ri:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lfd�uq ~ O   t cranstonw  Rsq ~ '1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_diego_cat san_diego_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~ Qq ~ �q ~ �t diegow  sq ~ 'n�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
des_moinest des_moines:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�|�Cuq ~ O   q ~�q ~�w  osq ~ '�e�esq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
atlanta_gat atlanta_ga:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�NI�uq ~ O   t atlantaw  �sq ~ '̤��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt west_valley_utt west_valley_ut:cxq ~q ~
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ Lޠe�uq ~ O   t westt valleyq ~�w  \sq ~ '�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt milwaukee_wit milwaukee_wi:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&sq ~ L�:�uq ~ O   t 	milwaukeet wiw  �sq ~ '��pq ~�sq ~ q ~q ~sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~0sq ~ L 3�uq ~ O   t manyw  	�sq ~ 'i���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt anderson_int anderson_in:cxq ~8q ~7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Asq ~ LǨ�uq ~ O   t andersonw  4sq ~ '7�8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt north_little_rock_art north_little_rock_ar:cxq ~Iq ~Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rsq ~ Li��Xuq ~ O   q ~ Qq ~ �t northq ~�q ~�w  bsq ~ 'K候sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt kalamazoo_mit kalamazoo_mi:cxq ~Zq ~Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~csq ~ L]���uq ~ O   q ~ Qq ~ �t 	kalamazoow  Csq ~ 'KH0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt schenectady_nyt schenectady_ny:cxq ~kq ~jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tsq ~ L���uq ~ O   t schenectadyw  @sq ~ 'w�u�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt troy_mit 	troy_mi:cxq ~|q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ln�uq ~ O   q ~ Qq ~ �t troyw  	Jsq ~ '9�ۑsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt hollywood_flt hollywood_fl:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LV��}uq ~ O   t 	hollywoodw  msq ~ '�qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt costa_mesa_cat costa_mesa_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LO�Duq ~ O   t costat mesaq ~"w  �sq ~ 'I/>�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	fresno_cat fresno_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��m�uq ~ O   t fresnow  Rsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	canton_oht canton_oh:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���'uq ~ O   q ~ Qq ~ �t cantonw  �sq ~ '�c�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt alhambra_cat alhambra_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lp�c�uq ~ O   q ~ Qq ~ �t alhambraw   msq ~ '�<��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
lansing_mit lansing_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L<�q�uq ~ O   t lansingq ~ gw  �sq ~ '0]��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t west_virginiat west_virginia:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LcZ�6uq ~ O   q ~t virginiaw  sq ~ '@��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt abingdon_pat abingdon_pa:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L����uq ~ O   t abingdonq ~w  �sq ~ 'n�zfsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t 	red_rivert red_river:rxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LA0Juq ~ O   q ~ Qt redq ~ �w   �sq ~ ';tn2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	nashua_nht nashua_nh:cxq ~'q ~&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0sq ~ L\)��uq ~ O   t nashuaq ~�t 	hampshirew  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt paterson_njt paterson_nj:cxq ~9q ~8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Bsq ~ L����uq ~ O   t patersonq ~�t jerseyw  �sq ~ '�w'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t kentuckyt 
kentucky:sxq ~Kq ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L�/��uq ~ O   q ~ Rq ~ Sq ~Mw  �sq ~ 'Q9sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t new_hampshiret new_hampshire:sxq ~[q ~Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ L��Kuq ~ O   q ~�q ~4w  8sq ~ '7���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt west_allis_wit west_allis_wi:cxq ~kq ~jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tsq ~ LvXhyuq ~ O   q ~t allist 	wisconsinw  �sq ~ '[A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt grand_prairie_txt grand_prairie_tx:cxq ~}q ~|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L׿�uq ~ O   q ~ Qq ~ �t grandt prairiew  (sq ~ '�L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
huntingtont huntington:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LU�W�uq ~ O   q ~�w  Usq ~ '�i�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5   lt lq ~ :q ~"t red:lxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L!\�uq ~ O   q ~q ~"w  �sq ~ 'sR��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t boiset boise:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Luq ~ O   q ~�w  	�sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt davenport_iat davenport_ia:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LhF'uq ~ O   q ~ Qq ~ �t 	davenportw  �sq ~ '�&{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt albuquerque_nmt albuquerque_nm:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��b�uq ~ O   t albuquerqueq ~�t mexicow  [sq ~ 'E�Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	newton_mat newton_ma:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lʹ�Wuq ~ O   q ~ Qq ~ �t newtonw  Osq ~ '`ْ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt santa_rosa_cat santa_rosa_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LD��uq ~ O   q ~ Qq ~ �t santat rosaw  �sq ~ '��-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt westminster_cat westminster_ca:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�\��uq ~ O   t westminsterq ~ �w  �sq ~ '� �7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~t pennsylvania:sxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L.���uq ~ O   q ~q ~ Rw   �sq ~ '9j �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt minneapolis_mnt minneapolis_mn:cxq ~&q ~%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/sq ~ L
�KSuq ~ O   t minneapolist 	minnesotaw  vsq ~ 'Þ\�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt great_falls_mtt great_falls_mt:cxq ~8q ~7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Asq ~ L6ٻ�uq ~ O   q ~ Qq ~ �t greatt fallsw  �sq ~ '%ڠ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	monroe_lat monroe_la:cxq ~Jq ~Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ssq ~ L�P'zuq ~ O   t monroew  �sq ~ '21;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t east_oranget east_orange:nxq ~[q ~Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ LɛE�uq ~ O   t eastt orangew  �sq ~ 'cM^q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~lq ~ksq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~psq ~ L�9 uq ~ O   t adjoinw  
Ksq ~ '��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~ysq ~ L�^�uq ~ O   q ~ �w  
,sq ~ '�w��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt irondequoit_nyt irondequoit_ny:cxq ~�q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L/�d1uq ~ O   q ~ Qq ~ �t irondequoitw  Ksq ~ 'M%��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt scottsdale_azt scottsdale_az:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�߲huq ~ O   t 
scottsdalew  �sq ~ '��J;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
hayward_cat hayward_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�ޢuq ~ O   t haywardq ~ �w  sq ~ '�U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
fremont_cat fremont_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   t fremontw  �sq ~ '+�T�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
alameda_cat alameda_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LY(��uq ~ O   t alamedaq ~ �w  	sq ~ 'xR�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t buffalot 	buffalo:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~�w  sq ~ '��ոsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt greensboro_nct greensboro_nc:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���Xuq ~ O   t 
greensborow  �sq ~ '�o^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt pasadena_txt pasadena_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��Quq ~ O   t pasadenat txw  �sq ~ '��t|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t green_rivert green_river:rxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L �uq ~ O   q ~ Qt greenw  �sq ~ '%�(�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	dallas_txt dallas_tx:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"sq ~ LU�ȕuq ~ O   t dallasq ~w  �sq ~ '��q;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
oakland_cat oakland_ca:cxq ~*q ~)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3sq ~ Lҕ.zuq ~ O   t oaklandq ~ �w  _sq ~ 't�Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fairfield_cat fairfield_ca:cxq ~;q ~:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Dsq ~ LA:uuq ~ O   t 	fairfieldq ~"w   �sq ~ 'Tּ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt tampa_flt 
tampa_fl:cxq ~Lq ~Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Usq ~ L�e�uq ~ O   t tampaw   usq ~ '�(��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
delaware:nxq ~]q ~\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~esq ~ L0��quq ~ O   q ~�w  �sq ~ '߉�Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt mesa_azt 	mesa_az:cxq ~lq ~ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~usq ~ L 3$uq ~ O   q ~�w  sq ~ 'Ya�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_haven_ctt new_haven_ct:cxq ~|q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L${�uq ~ O   q ~�t havent connecticutw  �sq ~ '���Vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lafayette_lat lafayette_la:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�KL�uq ~ O   t 	lafayettew  �sq ~ 'A�Vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t missouri_rivert missouri_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LW��Buq ~ O   q ~ Qt missouriq ~ �w  2sq ~ '  x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~ L   �uq ~ O   t aw   $sq ~ 'M���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
raleigh_nct raleigh_nc:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L:-�`uq ~ O   t raleighw   �sq ~ 'j���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt royal_oak_mit royal_oak_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�$�Xuq ~ O   t royalt oakq ~ gw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t rio_grande_rivert rio_grande_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�<�uq ~ O   q ~ Qt riot grandeq ~ �w  wsq ~ 'Ň}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t munciet muncie:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��{wuq ~ O   q ~�w  �sq ~ '�}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt columbia_mot columbia_mo:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L���uq ~ O   q ~Xt mow  ;sq ~ '�:�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t warwickt 	warwick:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LC	��uq ~ O   q ~w  �sq ~ '4H�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t westlandt 
westland:nxq ~$q ~#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-sq ~ L�S�Xuq ~ O   q ~&w  Wsq ~ 'QDuTsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~4q ~3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:sq ~ L��uq ~ O   q ~Dq ~Et mtw  sq ~ '�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_jose_cat san_jose_ca:cxq ~Bq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ksq ~ L��Euq ~ O   q ~ �t joseq ~ �w  �sq ~ '��~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t illinoist 
illinois:sxq ~Sq ~Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\sq ~ L�ctuq ~ O   q ~ Qq ~ Rq ~ Sq ~Uw  hsq ~ '22�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt overland_park_kst overland_park_ks:cxq ~cq ~bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lsq ~ L�(��uq ~ O   t overlandt parkw  �sq ~ '~;�q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~tq ~ssq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~xsq ~ L���uq ~ O   q ~ Rw  	�sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t nevadat nevada:sxq ~q ~~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LPi|wuq ~ O   q ~ Rq ~ Sq ~�w  ,sq ~ '�~��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t montanat 	montana:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LI�v*uq ~ O   q ~�w  �sq ~ '�l�:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L*J�luq ~ O   q ~ Qq ~ �q ~�q ~�w  _sq ~ 'RF��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t 
ohio_rivert ohio_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L jZNuq ~ O   q ~ Qt ohiow  �sq ~ '(v�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lynchburg_vat lynchburg_va:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L#�uq ~ O   t 	lynchburgw  �sq ~ '�\�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt elizabeth_njt elizabeth_nj:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�!@�uq ~ O   t 	elizabethw  �sq ~ '$��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Ѥ uq ~ O   q ~ Qq ~ Rq ~ Sq ~�q ~4w  �sq ~ '}�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt 
mount_yalet mount_yale:mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���huq ~ O   q ~ zt yalew  �sq ~ 'z�(4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_francisco_cat san_francisco_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	sq ~ L��vuq ~ O   q ~ �t 	franciscoq ~"w  �sq ~ '��
�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt penn_hills_pat penn_hills_pa:cxq ~	q ~	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	sq ~ L�.ϋuq ~ O   t pennt hillsq ~w  �sq ~ '�<2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ �I:�t 	<<e,t>,i>q ~ �q ~t countt count:<<e,t>,i>xq ~	 q ~	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   sq ~ �I:��t 	<<e,t>,e>q ~ �q ~ <xq ~	+sq ~ L!N�uq ~ O   t leastw   Rsq ~ '�y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t connecticut:sxq ~	5q ~	4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	=sq ~ Lf�1auq ~ O   q ~�w  Asq ~ '�s�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fall_river_mat fall_river_ma:cxq ~	Dq ~	Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	Msq ~ LC�uq ~ O   t fallq ~ �w  nsq ~ 'm~UJsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt redondo_beach_cat redondo_beach_ca:cxq ~	Uq ~	Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	^sq ~ L� �.uq ~ O   t redondot beachq ~"w  1sq ~ '+��Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt oak_lawn_ilt oak_lawn_il:cxq ~	gq ~	fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	psq ~ L{<!�uq ~ O   q ~ Qq ~ �q ~�t lawnw  csq ~ '�4K�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	newark_njt newark_nj:cxq ~	xq ~	wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ Lʹ]^uq ~ O   q ~ Qq ~ �t newarkw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bellevue_wat bellevue_wa:cxq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ Lau��uq ~ O   q ~�w  ksq ~ ':T��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt columbus_oht columbus_oh:cxq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ L��Quq ~ O   t columbust ohw  	sq ~ ',S�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~	�sq ~ L+ېuq ~ O   t locatedw  	�sq ~ 'x���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cambridge_mat cambridge_ma:cxq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ L��Vuq ~ O   t 	cambridgew  �sq ~ '��Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ LC�n�uq ~ O   q ~ Qq ~ �q ~�q ~�w  �sq ~ 'O���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	mobile_alt mobile_al:cxq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ L̃Fuq ~ O   q ~ Qq ~ �q ~w  _sq ~ '�P�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ Ldt�&uq ~ O   q ~�w  Asq ~ 'ĩ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 
new_mexicot new_mexico:sxq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~	�sq ~ L��2�uq ~ O   q ~�q ~�w  �sq ~ '$��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt corpus_christi_txt corpus_christi_tx:cxq ~	�q ~	�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
sq ~ Le��duq ~ O   t corpust christiw  "sq ~ '9ij[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt wilmington_det wilmington_de:cxq ~
q ~
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
sq ~ L�2�uq ~ O   t 
wilmingtont dew  �sq ~ 'ky��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lakewood_cat lakewood_ca:cxq ~
#q ~
"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
,sq ~ L��)\uq ~ O   t lakewoodq ~"w  ?sq ~ '	�Ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
salinas_cat salinas_ca:cxq ~
4q ~
3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
=sq ~ L{Nq�uq ~ O   q ~ Qq ~ �t salinasw  ~sq ~ ' �E�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt anchorage_akt anchorage_ak:cxq ~
Eq ~
Dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
Nsq ~ L�� uq ~ O   t 	anchoraget akw  �sq ~ '�~�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
sacramentot sacramento:nxq ~
Wq ~
Vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
`sq ~ LQ<H�uq ~ O   q ~
Yw  Xsq ~ 'ܡ�Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt greenwich_ctt greenwich_ct:cxq ~
gq ~
fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
psq ~ LS�x	uq ~ O   t 	greenwichq ~�w  �sq ~ '��[Esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	6xq ~
xq ~
wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
~sq ~ Ly%��uq ~ O   q ~�q ~ Rw  �sq ~ '!0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	laredo_txt laredo_tx:cxq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ L�[�uq ~ O   t laredoq ~ �w  �sq ~ 'ް��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
st_paul_mnt st_paul_mn:cxq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ L{�Auq ~ O   q ~ Qq ~ �q ~Nt paulw   �sq ~ '�0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ L�xffuq ~ O   q ~q ~ �w  sq ~ '�w��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
5xq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ LS�(Cuq ~ O   q ~
@q ~"w  Psq ~ '�w�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt waterbury_ctt waterbury_ct:cxq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ L���uq ~ O   t 	waterburyq ~�w  sq ~ '�H5;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t south_dakotat south_dakota:nxq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ Lz�L�uq ~ O   t southt dakotaw  �sq ~ 'c�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt north_charleston_sct north_charleston_sc:cxq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ L#�Juq ~ O   q ~Uq ~�w  �sq ~ '��?}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	las_vegast las_vegas:nxq ~
�q ~
�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
�sq ~ L���uq ~ O   q ~�q ~�w  �sq ~ '�MB�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt beaumont_txt beaumont_tx:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L� �%uq ~ O   t beaumontq ~w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ Lߢ�uq ~ O   q ~q ~
w  Qsq ~ '_Y:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_bedford_mat new_bedford_ma:cxq ~"q ~!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+sq ~ Lm6�Vuq ~ O   q ~ Qq ~ �q ~�t bedfordw  msq ~ 'p?hOsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	albany_gat albany_ga:cxq ~3q ~2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<sq ~ L��u�uq ~ O   q ~ Qq ~ �t albanyw  jsq ~ '�2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ �^��pt <<e,t>,<<e,i>,e>>q ~ �sq ~ �H��	t 	<<e,i>,e>sq ~ �|�t <e,i>q ~ <q ~q ~ <t argmaxt argmax:<<e,t>,<<e,i>,e>>xq ~Dq ~Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   sq ~ �W�i�t <<e,t>,<<e,e>,e>>q ~ �sq ~ �HgKt 	<<e,e>,e>q ~q ~ <xq ~Ssq ~ L�a�uq ~ O   t longestw   #sq ~ 'K+�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
bridgeportt bridgeport:nxq ~_q ~^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hsq ~ L�hO�uq ~ O   q ~aw  $sq ~ 'Ug�Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~oq ~nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~usq ~ L���_uq ~ O   q ~ Qq ~ �q ~�w  psq ~ '�v3Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~|q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�D<�uq ~ O   q ~ �q ~ Rw  $sq ~ '[OZsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t 
gila_rivert gila_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~ Qt gilaq ~ �w  �sq ~ '��zJq ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ ��%t <m,t>q ~ nq ~ �t mountaint mountain:<m,t>xq ~�q ~�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ L 4quq ~ O   t peakw  
Esq ~ '��,^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
danbury_ctt danbury_ct:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LU��)uq ~ O   t danburyw  �sq ~ '}��=q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~�q ~�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ L�%Cuq ~ O   t flowsw  	�sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	dayton_oht dayton_oh:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LVT�buq ~ O   t daytonq ~	�w  \sq ~ '!��6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	peoria_ilt peoria_il:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��9�uq ~ O   t peoriaw  �sq ~ 'c]'Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
detroit_mit detroit_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Li3_uq ~ O   q ~ Qq ~ �t detroitw  Rsq ~ 'Uagsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt kansas_city_kst kansas_city_ks:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�W�Muq ~ O   t kansasq ~ �q ~w  �sq ~ '�7H�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	cicero_ilt cicero_il:cxq ~
q ~	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�d)uq ~ O   q ~ Qq ~ �t cicerow  9sq ~ '�_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt elgin_ilt 
elgin_il:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$sq ~ L]>�Fuq ~ O   t elginq ~Uw  osq ~ '
�r{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~,q ~+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2sq ~ L-؎uq ~ O   q ~t ilw  �sq ~ ',�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~:q ~9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@sq ~ L\,�uq ~ O   q ~%q ~ �w  �sq ~ '�+-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
wyoming_mit wyoming_mi:cxq ~Gq ~Fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Psq ~ LBuq ~ O   t wyomingt miw  %sq ~ 'Bw�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~xt wisconsin:nxq ~Yq ~Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~asq ~ L��Suuq ~ O   q ~xw  #sq ~ '��E�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_britain_ctt new_britain_ct:cxq ~hq ~gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qsq ~ L�uq ~ O   q ~�t britaint ctw  �sq ~ '��l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_anterot mount_antero:mxq ~zq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ll�uq ~ O   q ~ zt anterow  �sq ~ ':�هsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LP�suq ~ O   q ~�q ~ �w  >sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~t utah:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�$��uq ~ O   q ~ Rq ~ Sq ~w  Gsq ~ '/P�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt st_joseph_mot st_joseph_mo:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lc���uq ~ O   q ~Nt josephq ~�w  3sq ~ '(���q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ �t majort major:<lo,t>xq ~�q ~�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ L }>uq ~ O   t bigw  
sq ~ 'E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~}xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��0Duq ~ O   q ~�q ~ gw  	�sq ~ '�Cdsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~Ft argmint argmin:<<e,t>,<<e,i>,e>>q ~	!xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~�sq ~ LW��uq ~ O   q ~ Qq ~	0w   Usq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t virginia_beacht virginia_beach:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L<���uq ~ O   q ~ q ~	bw  �sq ~ '�J�Vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t cimarron_rivert cimarron_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L0�rBuq ~ O   q ~ Qt cimarronq ~ �w  �sq ~ '�!jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
sq ~ L���uq ~ O   q ~w  �sq ~ '蓿\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t columbia_rivert columbia_river:rxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��quq ~ O   q ~ Qq ~Xw  �sq ~ '4^��q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ 8t floridat 	florida:sxq ~ q ~sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'sq ~ L 6M�uq ~ O   t thatw  
0sq ~ 'f��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bloomington_mnt bloomington_mn:cxq ~/q ~.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8sq ~ L�̵>uq ~ O   t bloomingtonq ~3w  5sq ~ 'c�5Nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ ��7��t 	<i,<i,t>>q ~sq ~ �}�t <i,t>q ~q ~ �t >t >:<i,<i,t>>sq ~ 0q ~t 	elevationt elevation:<lo,i>q ~Hxq ~@q ~?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~ �q ~q ~xq ~Psq ~ L6ǁ�uq ~ O   t highert thanw   Psq ~ '��Q(q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ Zt dover_det 
dover_de:cxq ~Xq ~Wsq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_sq ~ L�kvuq ~ O   t doverw  
4sq ~ '�\��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~gq ~fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~msq ~ Ly�/uq ~ O   q ~�t azw  2sq ~ ' ��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'xq ~uq ~tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{sq ~ L���"uq ~ O   q ~2t mnw   �sq ~ 'v���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt provo_utt 
provo_ut:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��m�uq ~ O   t provoq ~w  �sq ~ '�0ȅsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
abilene_txt abilene_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�q��uq ~ O   t abilenew  8sq ~ '��Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt tulsa_okt 
tulsa_ok:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��=uq ~ O   q ~ Qq ~ �t tulsaw  �sq ~ 'x��ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~ gt 
michigan:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�M�uq ~ O   q ~ gq ~ Rw  �sq ~ 'Cb�ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	winnebagot winnebago:lxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L	�z�uq ~ O   q ~q ~�w  �sq ~ 'AL4�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt brownsville_txt brownsville_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LM��uq ~ O   t brownsvilleq ~w  sq ~ 'X�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��dquq ~ O   q ~ Rq ~ Sq ~ �w  	sq ~ '�TՖsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~ Qq ~ �q ~	�w  jsq ~ '�_mYsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t 
missouri:sxq ~ q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LQy�uq ~ O   q ~�q ~ Rw  �sq ~ '���osq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t garden_grovet garden_grove:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�~Z�uq ~ O   t gardent grovew  �sq ~ '��I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t coloradot 
colorado:sxq ~!q ~ sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*sq ~ L5Z1Ruq ~ O   q ~ Qq ~ Rq ~ Sq ~#w  	�sq ~ '*;�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t santa_clarat santa_clara:nxq ~1q ~0sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:sq ~ L�m�zuq ~ O   q ~ t claraw  "sq ~ '�3��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt waterloo_iat waterloo_ia:cxq ~Bq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ksq ~ L �3uq ~ O   t waterloow  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t jacksont 	jackson:nxq ~Sq ~Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\sq ~ L���uq ~ O   q ~Uw  �sq ~ 'ևH�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
new_jerseyt new_jersey:nxq ~cq ~bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lsq ~ L���uq ~ O   q ~�q ~Fw  sq ~ 'o�ˠq ~�sq ~ q ~q ~sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~tsq ~ L��2�uq ~ O   t peoplew  	�sq ~ '���nq ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ ��Bt <p,t>sq ~ 5   pt pq ~ :q ~ �t placet place:<p,t>xq ~{q ~zsq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ L��.�uq ~ O   q ~Iw  	�sq ~ '���Bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt terre_haute_int terre_haute_in:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lb.nJuq ~ O   t terret hauteq ~w  �sq ~ '#W=4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt kansas_city_mot kansas_city_mo:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�3O�uq ~ O   q ~q ~ �w  sq ~ '760�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bridgeport_ctt bridgeport_ct:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L'��uq ~ O   q ~aq ~uw  �sq ~ '�E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	austin_txt austin_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�nh*uq ~ O   t austinq ~w  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LfH�uq ~ O   q ~t paw  �sq ~ '"�v�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt high_point_nct high_point_nc:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���tuq ~ O   t hight pointq ~Ut carolinaw  lsq ~ 'W�]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
Fxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L	�.�uq ~ O   q ~ Qq ~ �q ~
Qw  	sq ~ '-n8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t honolulut 
honolulu:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�Ruq ~ O   q ~ w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t hawaiit hawaii:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�z!uq ~ O   q ~w  	usq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	carson_cat carson_ca:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'sq ~ L�|=|uq ~ O   t carsonw  rsq ~ 'c�'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~/q ~.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5sq ~ L 6%�uq ~ O   q ~Nq ~
�w  vsq ~ '9ڗsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt southfield_mit southfield_mi:cxq ~<q ~;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Esq ~ L0,�uq ~ O   t 
southfieldw  �sq ~ 'ܵ*Dq ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ ���Dt 	<s,<c,t>>q ~ 8sq ~ �{6ot <c,t>q ~ Zq ~ �t capital2t capital2:<s,<c,t>>q ~�xq ~Lq ~Ksq ~ @q ~�sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~Wsq ~ L �Puq ~ O   q ~�w  
^sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
chicago_ilt chicago_il:cxq ~^q ~]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gsq ~ L-%Auq ~ O   t chicagoq ~Uw  vsq ~ '�C(�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
norwalk_cat norwalk_ca:cxq ~oq ~nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xsq ~ L�ܾuq ~ O   q ~ Qq ~ �t norwalkw  	�sq ~ '�&*Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt arlington_heights_ilt arlington_heights_il:cxq ~�q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L+@uq ~ O   t 	arlingtont heightsw  �sq ~ '�.ݛsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	aurora_ilt aurora_il:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�^)�uq ~ O   t auroraq ~5w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	taylor_mit taylor_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   t taylorq ~Tw   �sq ~ 'Iȩsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t snake_rivert snake_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Z�uq ~ O   q ~ Qt snakew  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~�sq ~ L6�0�uq ~ O   t highestw   Asq ~ 'L�4Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t parmat parma:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LX3uq ~ O   q ~�w  esq ~ '�L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�v�tuq ~ O   q ~ Qq ~ �q ~)w  `sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LG�J�uq ~ O   q ~w  		sq ~ 'u���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�uuq ~ O   q ~�q ~�w  �sq ~ 'U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
5xq ~
q ~	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ Ls�-�uq ~ O   q ~
@q ~ �w  	sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t lake_charlest lake_charles:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ sq ~ L2,�5uq ~ O   q ~t charlesw  �sq ~ '�_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt macon_gat 
macon_ga:cxq ~(q ~'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1sq ~ L-��uq ~ O   t maconw  esq ~ 't�7�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ �� t <r,t>q ~ �q ~ �q ~ �t river:<r,t>xq ~9q ~8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Csq ~ Lw�Juq ~ O   q ~ �w   ^sq ~ 'Q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~]t new_hampshire:nxq ~Jq ~Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rsq ~ L��Kuq ~ O   q ~�q ~4w  Bsq ~ '�_xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t seattlet 	seattle:nxq ~Yq ~Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bsq ~ LuSyuq ~ O   q ~[w  �sq ~ '�m�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt akron_oht 
akron_oh:cxq ~iq ~hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~rsq ~ L��y2uq ~ O   t akronq ~	�w  �sq ~ '��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t bakersfieldt bakersfield:nxq ~zq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�c��uq ~ O   q ~|w  �sq ~ '�"X�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
clifton_njt clifton_nj:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L?���uq ~ O   q ~ Qq ~ �t cliftonw  "sq ~ 'ک�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t bethesdat 
bethesda:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ln��`uq ~ O   q ~�w  �sq ~ 'يa�q ~Asq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ ���t <r,i>q ~ �q ~t lent 	len:<r,i>xq ~�q ~�sq ~ @q ~Osq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~�q ~Xw   5sq ~ '�Jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cedar_rapids_iat cedar_rapids_ia:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lv��Duq ~ O   t cedart rapidsw  4sq ~ 'w?�5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt sunnyvale_cat sunnyvale_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�<F�uq ~ O   t 	sunnyvaleq ~"w  sq ~ '�;��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt billings_mtt billings_mt:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LAH��uq ~ O   q ~ Qq ~ �t billingsw  $sq ~ 'ja�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fort_wayne_int fort_wayne_in:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�i[uq ~ O   q ~ �t waynew  sq ~ '����q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ ���t <t,t>q ~ �q ~ �t nott 	not:<t,t>xq ~�q ~�sq ~ @q ~�sq ~ G���    sq ~ sq ~ J   w   q ~�xq ~sq ~ L ��uq ~ O   t hasw  
Hsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�]uq ~ O   q ~ Qq ~Xq ~ �w  	ksq ~ 'yn+[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	odessa_txt odessa_tx:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#sq ~ L�=��uq ~ O   t odessaq ~w  'sq ~ '\v��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt koolaupoko_hit koolaupoko_hi:cxq ~+q ~*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4sq ~ LlMG�uq ~ O   t 
koolaupokow  csq ~ 'Gބ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~<q ~;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Bsq ~ LS��uq ~ O   q ~�q ~ �w  <sq ~ '��}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	euclid_oht euclid_oh:cxq ~Iq ~Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rsq ~ L�1H�uq ~ O   q ~ Qq ~ �t euclidw  �sq ~ 'ޣ�q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~t areat area:<lo,i>xq ~Yq ~Xsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~`sq ~ L -��uq ~ O   q ~[w  	�sq ~ 'NS�Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~gq ~fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~msq ~ LI0uq ~ O   q ~�q ~�w  	�sq ~ '��5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t upper_darbyt upper_darby:nxq ~tq ~ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}sq ~ LӴ�*uq ~ O   t uppert darbyw  �sq ~ '�>�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t rhode_islandt rhode_island:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LɠTuq ~ O   t rhodet islandq ~ Rw  Fsq ~ '��ĭsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt wichita_falls_txt wichita_falls_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lm�|~uq ~ O   t wichitaq ~Eq ~ �w  �sq ~ 'E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t massachusettst massachusetts:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��B�uq ~ O   q ~�w  fsq ~ '�޸Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t oklahomat 
oklahoma:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�x�uq ~ O   q ~�w  nsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L 6�Duq ~ O   q ~w  sq ~ 'P⾎sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fort_collins_cot fort_collins_co:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�>�Quq ~ O   q ~ Qq ~ �q ~ �t collinsw  dsq ~ 'b[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
garland_txt garland_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L �eguq ~ O   q ~ Qq ~ �t garlandw  	Usq ~ '
̧3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt columbia_sct columbia_sc:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L���uq ~ O   q ~ Qq ~ �q ~Xw  &sq ~ ' 19�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~sq ~ L 0��uq ~ O   t havew   sq ~ 'w���q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~q ~sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~sq ~ L ��uq ~ O   t liew  
Qsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t north_carolinat north_carolina:sxq ~!q ~ sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*sq ~ L�/uq ~ O   q ~Uq ~�w  �sq ~ '��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt mount_vernon_nyt mount_vernon_ny:cxq ~1q ~0sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:sq ~ L_		uq ~ O   q ~ zq ~�q ~�w  psq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t hartfordt 
hartford:nxq ~Aq ~@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ L��tuq ~ O   q ~Cw  �sq ~ '85$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt farmington_hills_mit farmington_hills_mi:cxq ~Qq ~Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Zsq ~ L�<�+uq ~ O   t 
farmingtonq ~	w  Qsq ~ '��B{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bakersfield_cat bakersfield_ca:cxq ~bq ~asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ksq ~ L�c��uq ~ O   q ~|w  �sq ~ '�(C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~rq ~qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xsq ~ L���uq ~ O   q ~�q ~�q ~�w   sq ~ 'l�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_blackburnt mount_blackburn:mxq ~q ~~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�5uq ~ O   q ~ zt 	blackburnw  -sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	kenner_lat kenner_la:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lȑ�kuq ~ O   q ~ Qq ~ �t kennerw  �sq ~ '�~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t whittiert 
whittier:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~�w  �sq ~ '�g �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t trentont 	trenton:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��X�uq ~ O   q ~�w  �sq ~ 'k��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lu� uq ~ O   q ~
�q ~uw  �sq ~ '��ϻsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�D�uq ~ O   q ~|q ~ �w  ,sq ~ 'P�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt sacramento_cat sacramento_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LQ<H�uq ~ O   q ~
Yw  �sq ~ '%]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t mississippit mississippi:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L߸�$uq ~ O   q ~�q ~ Rw  �sq ~ ' #Pq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~ L �uq ~ O   q ~ w  
Msq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~	sq ~ L�,Kuq ~ O   t withq ~ Qw   sq ~ ' dx.sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~sq ~ L c��uq ~ O   t howq ~3w    sq ~ '�s��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt utica_nyt 
utica_ny:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ L߀,uq ~ O   q ~ Qq ~ �t uticaw  >sq ~ '5��Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	downey_cat downey_ca:cxq ~0q ~/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9sq ~ L�1zuq ~ O   q ~ Qq ~ �t downeyw  tsq ~ '�+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
spokane_wat spokane_wa:cxq ~Aq ~@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ L�ٲ}uq ~ O   t spokanew  	sq ~ '�X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fayetteville_nct fayetteville_nc:cxq ~Rq ~Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[sq ~ L�̩�uq ~ O   t fayettevillet ncw  gsq ~ '0��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt charlotte_nct charlotte_nc:cxq ~dq ~csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~msq ~ L]�[)uq ~ O   t 	charlotteq ~_w  �sq ~ 'm�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~uq ~tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{sq ~ L@��iuq ~ O   q ~�q ~ gw  �sq ~ '�)'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	eugene_ort eugene_or:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   t eugenew  sq ~ '|��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t philadelphiat philadelphia:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LR`6suq ~ O   q ~�w  �sq ~ '�,h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
compton_cat compton_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L8��"uq ~ O   t comptonw  Usq ~ '���asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~jxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��tuq ~ O   q ~uq ~�w  	sq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt niagara_falls_nyt niagara_falls_ny:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��P�uq ~ O   t niagaraq ~Eq ~�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lu��uq ~ O   q ~ q ~q ~ �w  sq ~ ')=pHsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L[&�uq ~ O   q ~Uq ~�q ~�q ~fw  �sq ~ '�p#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~qw  wsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt irvington_njt irvington_nj:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L-�Yuq ~ O   t 	irvingtonw  #sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<xq ~
q ~	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�[��uq ~ O   q ~Gw  ;sq ~ '�۠[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�G8�uq ~ O   q ~Nt iaw  Lsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lynn_mat 	lynn_ma:cxq ~%q ~$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.sq ~ Ló�uq ~ O   t lynnq ~�w  Xsq ~ '�s��q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~5q ~4sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~9sq ~ LL�E�uq ~ O   t traversew  
[sq ~ '�<.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t arkansas_rivert arkansas_river:rxq ~Aq ~@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ L�/�uq ~ O   q ~ Qq ~fw  �sq ~ '�G9q ~�sq ~ sq ~ sq ~ J   w   q ~Eq ~�xq ~Pq ~Osq ~ @q ~�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~Tsq ~ L��auq ~ O   t unitedw  
sq ~ ' �Mq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~]sq ~ L �uq ~ O   t canw  	�sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t idahot idaho:sxq ~eq ~dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~nsq ~ L��kuq ~ O   q ~gw  �sq ~ '�4 sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt appleton_wit appleton_wi:cxq ~uq ~tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~sq ~ L}~uq ~ O   t appletonq ~xw  �sq ~ 'i�$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 
washingtont washington:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��yuq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  	Rsq ~ '(I�}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t smoky_hill_rivert smoky_hill_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�6!�uq ~ O   q ~ Qt smokyt hillw  �sq ~ 'Io�ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt westland_mit westland_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LM�Ruq ~ O   q ~&q ~ gw   �sq ~ '���Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
redford_mit redford_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L@�
uq ~ O   t redfordw  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt greenville_sct greenville_sc:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�O��uq ~ O   q ~ Qq ~ �t 
greenvillew  tsq ~ '^�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	lexingtont lexington:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Nuq ~ O   q ~�w  :sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
hampton_vat hampton_va:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L[��nuq ~ O   t hamptonq ~ w  rsq ~ '�U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~5t tennessee:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LGdg]uq ~ O   q ~5q ~ Rw  �sq ~ '~B��q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~	q ~sq ~ @q ~ �sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~q ~ �w   sq ~ 'vk�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ Lř�uq ~ O   q ~�q ~�w   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt huntington_beach_cat huntington_beach_ca:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ L��̷uq ~ O   q ~�q ~	bq ~"w  �sq ~ '��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt santa_monica_cat santa_monica_ca:cxq ~/q ~.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8sq ~ L���Nuq ~ O   q ~ t monicaq ~ �w  �sq ~ '��i[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt huntsville_alt huntsville_al:cxq ~@q ~?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Isq ~ L|�>9uq ~ O   t 
huntsvillet alw  tsq ~ '|
4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t jacksonvillet jacksonville:nxq ~Rq ~Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[sq ~ Lg�zuq ~ O   q ~Tw   �sq ~ 'p*�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt scotts_valley_cat scotts_valley_ca:cxq ~bq ~asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ksq ~ L����uq ~ O   t scottsq ~q ~ �w  !sq ~ '�e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~xt wisconsin:sxq ~sq ~rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{sq ~ L��Yuq ~ O   q ~ Rq ~ Sq ~xw  zsq ~ '㨷�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
houston_txt houston_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LA�Ōuq ~ O   t houstonw   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�A�uq ~ O   q ~3w  	Csq ~ '�p��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt stamford_ctt stamford_ct:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lw�|�uq ~ O   t stamfordq ~uw  5sq ~ 'Ƥsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L|T��uq ~ O   q ~	q ~	q ~�w  psq ~ '�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	norman_okt norman_ok:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L~���uq ~ O   q ~�t okw  �sq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	raleigh:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L:-�`uq ~ O   q ~�w  �sq ~ '�@�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~ L�@(uq ~ O   t pleasew   	sq ~ 'AY7�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t renot reno:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L 5[ruq ~ O   q ~�w  �sq ~ '�n�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt little_rock_art little_rock_ar:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LXo�`uq ~ O   q ~�q ~�q ~ �w  �sq ~ '�  �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~
�t south_dakota:sxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��uq ~ O   q ~
�q ~
�q ~ Rw  sq ~ '��v;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t north_dakotat north_dakota:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$sq ~ Lr4�Iuq ~ O   q ~Uq ~
�w  Isq ~ 'ۏ`>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t west_virginia:sxq ~+q ~*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3sq ~ L��yuq ~ O   q ~q ~ q ~ Rw  Msq ~ ''	�0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt springfield_ilt springfield_il:cxq ~:q ~9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Csq ~ L�1�Kuq ~ O   t springfieldw  1sq ~ '�'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt oceanside_cat oceanside_ca:cxq ~Kq ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L _�uq ~ O   t 	oceansidew  �sq ~ '�Z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt gary_int 	gary_in:cxq ~\q ~[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~esq ~ Ly��uq ~ O   t garyt indianaw   �sq ~ 'H�k:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~nq ~msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tsq ~ L���uq ~ O   q ~ Qq ~ �q ~q ~ww  Msq ~ 'd��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t nebraskat 
nebraska:nxq ~{q ~zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L/E�uq ~ O   q ~}w   �sq ~ '�#�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t midlandt 	midland:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L>��quq ~ O   q ~�w  �sq ~ '^�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Nt 
waterloo:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L �3uq ~ O   q ~Nw  �sq ~ '�<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�eJuq ~ O   q ~ Qq ~ �q ~�w  msq ~ '�a�Fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�3 iuq ~ O   q ~ Qq ~ �q ~�w  ~sq ~ '�#e+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t farmington_hillst farmington_hills:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�<�+uq ~ O   q ~]q ~	w  �sq ~ '
V,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_browne_towert mount_browne_tower:mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LY�Quq ~ O   q ~ zt brownet towerw  "sq ~ '&"Dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
kendall_flt kendall_fl:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LW/�uq ~ O   t kendallt flw  !sq ~ '�=Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t oregont oregon:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��ޢuq ~ O   q ~�w  Nsq ~ '��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	hxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ Lj*�uq ~ O   q ~�q ~	sq ~5w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t kansas_cityt kansas_city:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�3O�uq ~ O   q ~q ~ �w  sq ~ 'X4OJsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt st_petersburg_flt st_petersburg_fl:cxq ~%q ~$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.sq ~ L��(uq ~ O   q ~ Qq ~ �q ~Nq ~Ow  �sq ~ '�]�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lakewood_cot lakewood_co:cxq ~5q ~4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>sq ~ L��/uq ~ O   q ~
/t cow  vsq ~ '$�Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~t kansas:sxq ~Fq ~Esq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Nsq ~ LK4�uq ~ O   q ~ Rq ~ Sq ~w  sq ~ 'xr�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Vsq ~ Lw�Juq ~ O   q ~ �w  
sq ~ '�[Șsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	danbury:nxq ~]q ~\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~esq ~ LU��)uq ~ O   q ~�w  	sq ~ '��H�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~lq ~ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~rsq ~ LB�/�uq ~ O   q ~�q ~�q ~Uw  �sq ~ '��isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~yq ~xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L?u)uq ~ O   q ~Nq ~
�q ~3w  ksq ~ '�F�4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt baton_rouge_lat baton_rouge_la:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L3�Quq ~ O   t batont rouget 	louisianaw  �sq ~ '�~��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lake_charles_lat lake_charles_la:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L2,�5uq ~ O   q ~q ~#w  �sq ~ 'XWd|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�bDuq ~ O   q ~ Qq ~ �w  �sq ~ '��uXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	clifton:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L3L�uq ~ O   q ~�w  sq ~ 'G̽�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ls�~�uq ~ O   q ~ Rq ~ Sq ~�w  �sq ~ 'p�j|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t delaware_rivert delaware_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L0��uq ~ O   q ~ Qq ~�w  �sq ~ '1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~exq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L]�4*uq ~ O   q ~pw  rsq ~ 'i���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Dt 
anderson:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LǨ�uq ~ O   q ~Dw  [sq ~ '��<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t cheyenne_rivert cheyenne_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L]�uq ~ O   q ~ Qt cheyennew  �sq ~ 'Q<�
q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~sq ~ LQ<H�uq ~ O   q ~
Yw  
Bsq ~ '�x�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t colorado_rivert colorado_river:rxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ sq ~ Lڻ;�uq ~ O   q ~ Qq ~#w  4sq ~ '/9�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt newport_beach_cat newport_beach_ca:cxq ~'q ~&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0sq ~ L����uq ~ O   t newportq ~	bq ~ �w  �sq ~ '$ڕ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt hamilton_oht hamilton_oh:cxq ~8q ~7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Asq ~ L��gzuq ~ O   t hamiltonw  Csq ~ '�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
shreveportt shreveport:nxq ~Iq ~Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rsq ~ L��6uq ~ O   q ~Kw  &sq ~ '�l��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5  lt coq ~ :t usat usa:coxq ~Yq ~Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ L�Tuq ~ O   t continentalt usw  �sq ~ '���)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fullerton_cat fullerton_ca:cxq ~mq ~lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vsq ~ L�^��uq ~ O   t 	fullertonw  Jsq ~ '�$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	hayward:nxq ~~q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L)��Zuq ~ O   q ~�w  �sq ~ 'A��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t edisont edison:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~�w  sq ~ '�g�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�i�uq ~ O   q ~�q ~�q ~fw  Osq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��$uq ~ O   q ~ Qq ~ �q ~�q ~ �w  �sq ~ 'q�[5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t citrus_heightst citrus_heights:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L^��Juq ~ O   t citrusq ~�w  ysq ~ 'r$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ut 
illinois:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~Uw  �sq ~ '�BW�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
concord_cat concord_ca:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Dtuq ~ O   t concordq ~ �w  Usq ~ 'MoXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t bouldert 	boulder:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L/�+uq ~ O   q ~�w  �sq ~ '�Ƨisq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lexington_kyt lexington_ky:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��]�uq ~ O   q ~�q ~Mw  sq ~ '��rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt jacksonville_flt jacksonville_fl:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L]�^�uq ~ O   q ~Tq ~"w  �sq ~ 'ŘH@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt santa_ana_cat santa_ana_ca:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!sq ~ LD�auq ~ O   q ~ Qq ~ �q ~ t anaw  {sq ~ '��V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt santa_barbara_cat santa_barbara_ca:cxq ~)q ~(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2sq ~ L��U"uq ~ O   q ~ t barbaraq ~"w  Psq ~ '�q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	casper_wyt casper_wy:cxq ~:q ~9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Csq ~ L��GZuq ~ O   t casperq ~Sw  �sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt amarillo_txt amarillo_tx:cxq ~Kq ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L���guq ~ O   q ~ Qq ~ �t amarillow  ;sq ~ '�"Osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~\q ~[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bsq ~ L��w-uq ~ O   q ~Nq ~Oq ~"w  �sq ~ '2��~q ~�sq ~ sq ~ sq ~ J   w   q ~Hxq ~hq ~gsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~lsq ~ L��.�uq ~ O   q ~Iw  
sq ~ 'r7�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~sq ~rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ysq ~ L���uq ~ O   q ~Uw  	\sq ~ '1h��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt framingham_mat framingham_ma:cxq ~�q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��kJuq ~ O   t 
framinghamt maw  7sq ~ '��Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_brosst mount_bross:mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��˦uq ~ O   q ~ zt brossw  �sq ~ '�Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L/��uq ~ O   q ~�q ~pw  �sq ~ '�2��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��,uq ~ O   q ~�q ~�q ~ �w  �sq ~ '��)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t wateree_catawba_rivert wateree_catawba_river:rxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���Vuq ~ O   t watereet catawbaq ~ �w  �sq ~ '�ŭ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt worcester_mat worcester_ma:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L3���uq ~ O   t 	worcesterw  	Wsq ~ '��vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t venturat 	ventura:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�`�uq ~ O   q ~�w  (sq ~ '�� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt plano_txt 
plano_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�K
uq ~ O   q ~ Qq ~ �t planow  ;sq ~ '�9?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt upper_darby_pat upper_darby_pa:cxq ~q ~ sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
sq ~ L��euq ~ O   q ~�q ~�q ~�w  �sq ~ 'S�Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LGQ��uq ~ O   q ~5q ~ �w  �sq ~ '>rߵsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t neosho_rivert neosho_river:rxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'sq ~ Lt�
uq ~ O   t neoshoq ~ �w  sq ~ 'w�h]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~/q ~.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~5sq ~ L  cuq ~ O   q ~w   Dsq ~ '8���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt birmingham_alt birmingham_al:cxq ~<q ~;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Esq ~ L��Uuq ~ O   t 
birminghamt alabamaw  �sq ~ '\c�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Nq ~Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L�/��uq ~ O   q ~ Qq ~ �q ~�q ~Ew  sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt los_angeles_cat los_angeles_ca:cxq ~[q ~Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ L��uq ~ O   q ~/q ~0q ~"w  >sq ~ 'I� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t arlington:nxq ~kq ~jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ssq ~ Lz���uq ~ O   q ~�w  	+sq ~ 'SRI�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt pensacola_flt pensacola_fl:cxq ~zq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LB�5uq ~ O   t 	pensacolaq ~"w  �sq ~ '�۬�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	aurora_cot aurora_co:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�^(�uq ~ O   q ~�q ~Aw  �sq ~ '�|�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�I-uq ~ O   q ~�t iowaw  <sq ~ ' ��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~ L �Puq ~ O   q ~�w  
Ysq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
wichita_kst wichita_ks:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~�t ksw  �sq ~ '�Ӕ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t longviewt 
longview:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�jc_uq ~ O   q ~�w  7sq ~ '�S=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t grand_rapidst grand_rapids:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L~KCKuq ~ O   q ~�q ~�w  �sq ~ '�r*�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt tallahassee_flt tallahassee_fl:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�DX�uq ~ O   t tallahasseeq ~"w  �sq ~ '{9{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt tyler_txt 
tyler_tx:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���puq ~ O   t tylerq ~w   sq ~ 'qڐsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~
sq ~ LU�Xuq ~ O   q ~ q ~q ~"w  �sq ~ '�V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~sq ~ L���uq ~ O   t shortestw   sq ~ '9�	;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt columbus_gat columbus_ga:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ L��Ruq ~ O   q ~	�t gaw  !sq ~ '!.��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t roanoke_rivert roanoke_river:rxq ~0q ~/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9sq ~ L����uq ~ O   q ~ Qt roanokeq ~ �w  	sq ~ '<Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Aq ~@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Gsq ~ L(mSFuq ~ O   q ~�q ~Uq ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\xq ~Nq ~Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L���uq ~ O   q ~/q ~0q ~ �w  sq ~ '���q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~\sq ~ L��uq ~ O   t urbanw  
=sq ~ '@ik'q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ nt guadalupe_peakt guadalupe_peak:mxq ~cq ~bsq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jsq ~ L 4quq ~ O   q ~�w  
sq ~ '<T'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~qq ~psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wsq ~ L���uq ~ O   q ~ Qq ~ �q ~q ~#w  sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~~q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lqq�uq ~ O   q ~q ~uw  Wsq ~ '�'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t loraint lorain:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~�w  �sq ~ '+�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt hartford_ctt hartford_ct:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�i>�uq ~ O   q ~Cq ~uw  @sq ~ ']�}q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~�q ~�sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lm\4�uq ~ O   t 
kilometersw  
Ssq ~ '���Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~ Qq ~ Rq ~ Sq ~�q ~�w  	*sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	arvada_cot arvada_co:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��IPuq ~ O   t arvadaq ~#w  Zsq ~ 'B�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
orlando_flt orlando_fl:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L)WD�uq ~ O   t orlandoq ~"w  �sq ~ '5Jy�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t dulutht duluth:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�H:uq ~ O   q ~�w  �sq ~ '&�Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt arlington_vat arlington_va:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Q��uq ~ O   q ~�q ~=w  	?sq ~ '	�L�q ~�sq ~ sq ~ sq ~ J   w   q ~Eq ~xq ~q ~sq ~ @q ~�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~sq ~ L 3;�uq ~ O   t mostw  	�sq ~ '�j8xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t aurora:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�,S�uq ~ O   q ~�w  �sq ~ '�`J8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t austin:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'sq ~ L�,ٸuq ~ O   q ~�w  +sq ~ '��C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~.q ~-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4sq ~ LQ�8.uq ~ O   q ~ Qq ~<w  �sq ~ 'Pߋ�q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~Pt capitalt capital:<c,t>xq ~:q ~9sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Asq ~ L��uq ~ O   t largestw  
sq ~ '��4Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt sioux_city_iat sioux_city_ia:cxq ~Iq ~Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rsq ~ L����uq ~ O   t siouxq ~ �q ~ w  Gsq ~ 'Xb98sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~St 	wyoming:nxq ~Zq ~Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bsq ~ Lk�C�uq ~ O   q ~Sw  �sq ~ 'ǥ\q ~=sq ~ sq ~ sq ~ 
w   q ~Axq ~hq ~gsq ~ @q ~Lsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~lq ~Qw   ,sq ~ '99sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~qq ~psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wsq ~ L�r�Xuq ~ O   q ~Wq ~ Sq ~Xq ~ Rw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~~q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�=�uq ~ O   q ~Uq ~�q ~
�q ~�w  
sq ~ '�';sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
seattle_wat seattle_wa:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L5��uq ~ O   q ~[t waw  sq ~ '��Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt montgomery_alt montgomery_al:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�PLSuq ~ O   q ~ Qq ~ �t 
montgomeryw  6sq ~ 'Fݘsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t taylor:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lˁ�auq ~ O   q ~�w  sq ~ '��V2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt miami_flt 
miami_fl:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�N:<uq ~ O   t miamiq ~"w  	Gsq ~ '�O[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LI��uq ~ O   q ~q ~Mw  �sq ~ '~nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ L��%uq ~ O   t wherew   sq ~ '0U3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt champaign_ilt champaign_il:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LU��uq ~ O   t 	champaignw  ssq ~ 'M0�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ft kalamazoo:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LQ�k�uq ~ O   q ~fw  �sq ~ 'xHsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt east_los_angeles_cat east_los_angeles_ca:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L~�Zuq ~ O   q ~gq ~/q ~0w  ysq ~ '`�'2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt dearborn_heights_mit dearborn_heights_mi:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!sq ~ Ld�]uq ~ O   q ~ Qq ~ �q ~ fq ~�w  sq ~ '׫~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~t densityt density:<lo,i>xq ~(q ~'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~1sq ~ L��uq ~ O   q ~q ~*w   Wsq ~ '�=G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt allentown_pat allentown_pa:cxq ~8q ~7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Asq ~ L�h@uq ~ O   q ~ Qq ~ �t 	allentownw  �sq ~ 'rU��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
�t waterbury:nxq ~Iq ~Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Qsq ~ L�B��uq ~ O   q ~
�w  �sq ~ '�f)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Xq ~Wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^sq ~ L�b��uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��n�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t independencet independence:nxq ~eq ~dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~nsq ~ L �vZuq ~ O   q ~gw  `sq ~ '�[q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~vsq ~ L���uq ~ O   t whosew  	�sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~#t north_carolina:nxq ~~q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�/uq ~ O   q ~Uq ~�w  �sq ~ '��#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~�w   jsq ~ '��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt sterling_heights_mit sterling_heights_mi:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L� ��uq ~ O   t sterlingq ~�w  	osq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�!/Kuq ~ O   q ~w  �sq ~ ':	��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt virginia_beach_vat virginia_beach_va:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L<���uq ~ O   q ~ q ~	bw  sq ~ 'ڬ!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t berkeleyt 
berkeley:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lk�c�uq ~ O   q ~�w  Hsq ~ '���q ~�sq ~ sq ~ sq ~ J   w   q ~	!xq ~�q ~�sq ~ @q ~�sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�sq ~ L��3uq ~ O   q ~?w  
Osq ~ '��9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt rochester_nyt rochester_ny:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ln�I:uq ~ O   t 	rochesterq ~�w  	�sq ~ 'HSCsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bethesda_mdt bethesda_md:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L{X�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ 'gD��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt st_clair_shores_mit st_clair_shores_mi:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��6Vuq ~ O   q ~Nt clairt shoresq ~Tw  asq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	edison_njt edison_nj:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LU��uq ~ O   q ~�q ~�q ~Fw  �sq ~ 't�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~%q ~$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+sq ~ L�ҷuq ~ O   q ~4t georgiaw   �sq ~ 'c���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	tacoma_wat tacoma_wa:cxq ~3q ~2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<sq ~ L�w�+uq ~ O   t tacomaw  	Zsq ~ 'W��Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Dq ~Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ L�&Ouq ~ O   q ~�q ~�q ~iw  	Fsq ~ '�E�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Qq ~Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Wsq ~ LS��uq ~ O   q ~ Qq ~ �q ~w  �sq ~ '�r�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~it 	indiana:sxq ~^q ~]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fsq ~ L��uq ~ O   q ~ Rq ~ Sq ~iw  �sq ~ '�5>�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~mq ~lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ssq ~ L���.uq ~ O   q ~ Qq ~ �q ~aw  �sq ~ '���+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt knoxville_tnt knoxville_tn:cxq ~zq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L^��uq ~ O   t 	knoxvillew  ysq ~ 'W�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	quincy_mat quincy_ma:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LӮ1#uq ~ O   q ~ Qq ~ �t quincyw  �sq ~ '�6�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
phoenix_azt phoenix_az:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�8�juq ~ O   t phoenixq ~pw  �sq ~ '1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cincinnati_oht cincinnati_oh:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��7uq ~ O   t 
cincinnatiq ~�w  �sq ~ '�<�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��L�uq ~ O   q ~ �q ~w  �sq ~ '�}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	baltimoret baltimore:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L;���uq ~ O   q ~�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t new_yorkt 
new_york:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�D�uq ~ O   q ~�q ~�q ~ Rw  �sq ~ '4��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LJ�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�FЛsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_maroont mount_maroon:mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��Wuq ~ O   q ~ zt maroonw  �sq ~ 'l���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt st_louis_mot st_louis_mo:cxq ~	q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L����uq ~ O   q ~ Qq ~ �q ~Nt louisw  �sq ~ '�"l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Eq ~Hxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~ sq ~ L6�0�uq ~ O   q ~�w   ]sq ~ 'l���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~'q ~&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-sq ~ Lc��?uq ~ O   q ~�q ~	bw  �sq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~t sizet size:<lo,i>xq ~4q ~3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~=sq ~ L��uq ~ O   q ~Dw   Esq ~ '��<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt miami_beach_flt miami_beach_fl:cxq ~Dq ~Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Msq ~ L�^�uq ~ O   q ~�q ~	bq ~�w  �sq ~ '��dTsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Tq ~Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Zsq ~ L�5t.uq ~ O   q ~Nq ~�w  �sq ~ '��4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt shreveport_lat shreveport_la:cxq ~aq ~`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jsq ~ L��6uq ~ O   q ~Kw  �sq ~ ')u�qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~qq ~psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wsq ~ L�S�Xuq ~ O   q ~&w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~bxq ~~q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�>m�uq ~ O   q ~ Qq ~ �q ~Kw  5sq ~ '�.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t vermontt 	vermont:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Loǿ�uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  Nsq ~ '��|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ln
T!uq ~ O   q ~�q ~�w  �sq ~ 'YN��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t racinet racine:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~�w  Hsq ~ 'I�U[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t mountain_viewt mountain_view:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L{u�uq ~ O   q ~�t vieww  �sq ~ '�Bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L'W��uq ~ O   q ~ Qq ~ �q ~ �q ~ �w  �sq ~ 'M��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~_xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Ls��huq ~ O   q ~iw   psq ~ '�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	!xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�sq ~ L�8muq ~ O   t atq ~	0t onew   sq ~ 'XJsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���ruq ~ O   q ~Uq ~�q ~�w  nsq ~ '�ϱYsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ sq ~ L6'E�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ ',��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~ q ~ sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ sq ~ Lyp�$uq ~ O   q ~Nq ~q ~w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~ q ~ sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ sq ~ L��uq ~ O   q ~ Qq ~ �q ~	�w  sq ~ '�2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~ &q ~ %sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ ,sq ~ L���6uq ~ O   q ~ �q ~ �w  �sq ~ '闃xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ft casper:nxq ~ 3q ~ 2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ ;sq ~ L�|�fuq ~ O   q ~Fw  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt salem_ort 
salem_or:cxq ~ Bq ~ Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ Ksq ~ L���}uq ~ O   t salemq ~`w  psq ~ '���nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt santa_clara_cat santa_clara_ca:cxq ~ Sq ~ Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ \sq ~ L�h��uq ~ O   q ~ q ~=q ~"w  �sq ~ 'ջ:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~ cq ~ bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ isq ~ L�sóuq ~ O   q ~�w  	Ssq ~ 'æ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~ pq ~ osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ vsq ~ Lբpuq ~ O   q ~q ~w  )sq ~ '{�Xusq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~ }q ~ |sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L�+=Fuq ~ O   q ~Uq ~ Rw  �sq ~ 'H!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	Vxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ Lפ�uq ~ O   q ~	aq ~	bw  �sq ~ 'C���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	elyria_oht elyria_oh:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L��Y�uq ~ O   t elyriaq ~	�w  sq ~ '��&�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t burbankt 	burbank:nxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L>-yuq ~ O   q ~ �w  <sq ~ '�w��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
madison_wit madison_wi:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L����uq ~ O   t madisonq ~*w  �sq ~ '��	sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L{=>�uq ~ O   q ~ Qq ~ �q ~ �q ~Nw  	�sq ~ '�,W�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	royal_oakt royal_oak:nxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L��Ғuq ~ O   q ~�q ~�w  isq ~ '�[icsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t fort_collinst fort_collins:nxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L>i�uq ~ O   q ~ �q ~�w  ]sq ~ '��Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_orleans_lat new_orleans_la:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L3��duq ~ O   q ~ Qq ~ �q ~�t orleansw  �sq ~ '2+�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t sioux_fallst sioux_falls:nxq ~!q ~!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!sq ~ L�J|uq ~ O   q ~Uq ~Ew  �sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t wichita_fallst wichita_falls:nxq ~!q ~!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~! sq ~ L���uq ~ O   q ~�q ~Ew  Fsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
somervillet somerville:nxq ~!'q ~!&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!0sq ~ L�Ruq ~ O   q ~!)w  �sq ~ '~k;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_williamsont mount_williamson:mxq ~!7q ~!6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!@sq ~ L�_`Vuq ~ O   q ~ zt 
williamsonw  sq ~ 'B锲sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~ft 
arkansas:sxq ~!Hq ~!Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!Psq ~ L5�Vuq ~ O   q ~ Rq ~ Sq ~fw  sq ~ '"N�Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~!Wq ~!Vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!]sq ~ LMB��uq ~ O   q ~�q ~�w  2sq ~ '�9r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	muncie_int muncie_in:cxq ~!dq ~!csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!msq ~ L����uq ~ O   q ~�q ~iw  �sq ~ '5��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_leandro_cat san_leandro_ca:cxq ~!tq ~!ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!}sq ~ LD<i�uq ~ O   q ~ �t leandroq ~"w  �sq ~ '=�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ L|�$uq ~ O   q ~q ~wq ~*w  `sq ~ '  �\q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~!�sq ~ L  uq ~ O   t onw  	�sq ~ 'g�h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt port_arthur_txt port_arthur_tx:cxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ L�ɛ�uq ~ O   t portt arthurq ~w  	'sq ~ '�fv7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ L�M��uq ~ O   q ~ Qq ~Wt statesw  �sq ~ 'C�(8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t torrancet 
torrance:nxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ L�ضuq ~ O   q ~!�w  �sq ~ 'G�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
reading_pat reading_pa:cxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ L�T�uq ~ O   t readingq ~�w  	�sq ~ '�-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
saginaw_mit saginaw_mi:cxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ Lnϋ�uq ~ O   t saginaww  Bsq ~ ' �y�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt longview_txt longview_tx:cxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~!�sq ~ L����uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
bayonne_njt bayonne_nj:cxq ~!�q ~!�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"sq ~ L�܈>uq ~ O   t bayonneq ~�q ~Fw  sq ~ '�)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt clearwater_flt clearwater_fl:cxq ~"q ~"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"sq ~ L��g�uq ~ O   q ~ Qq ~ �t 
clearwaterw  1sq ~ '�`|�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~}xq ~"q ~"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"%sq ~ L��uq ~ O   q ~ Qq ~ �q ~�q ~�w  	=sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
norwalk_ctt norwalk_ct:cxq ~",q ~"+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"5sq ~ L[�'wuq ~ O   q ~{q ~uw  �sq ~ 'rL��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
ventura_cat ventura_ca:cxq ~"<q ~";sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"Esq ~ L�`�uq ~ O   q ~�w   �sq ~ '|�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t skokiet skokie:nxq ~"Lq ~"Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"Usq ~ L�U6�uq ~ O   q ~"Nw  8sq ~ '!�-q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~"]sq ~ L!���uq ~ O   t neighboringw  	�sq ~ '3��q ~�sq ~ sq ~ sq ~ J   w   q ~Msq ~ 0q ~ Zt 	albany_nyt albany_ny:cxq ~"dq ~"csq ~ @q ~�sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~"ksq ~ LL�E�uq ~ O   q ~<w  
Nsq ~ '���msq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
boulder_cot boulder_co:cxq ~"rq ~"qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"{sq ~ Lhf�uq ~ O   q ~ Qq ~ �q ~�w  isq ~ 'N�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t 
pasadena:nxq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ LG�J�uq ~ O   q ~w  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~bxq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ L�&��uq ~ O   q ~Kq ~�w  �sq ~ '>�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ L.� 3uq ~ O   q ~<w  �sq ~ '��%�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ Lp�>uq ~ O   q ~q ~#t law   |sq ~ '�x�$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t lake_of_the_woodst lake_of_the_woods:lxq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ L��,
uq ~ O   q ~q ~q ~ Sq ~ Qt woodsw  	�sq ~ '��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~"�sq ~ Lї�uq ~ O   t foundw  
sq ~ '�7�Asq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lakewood_oht lakewood_oh:cxq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ L��+cuq ~ O   q ~
/q ~�w  �sq ~ '�ի�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t potomac_rivert potomac_river:rxq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ L;��uq ~ O   q ~ Qt potomacq ~ �w  �sq ~ '� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2xq ~"�q ~"�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"�sq ~ L����uq ~ O   q ~ zq ~�q ~�q ~�w  �sq ~ '��?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t camdent camden:nxq ~#q ~# sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#
sq ~ L�y�uq ~ O   q ~#w  sq ~ '킯�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	green_bayt green_bay:nxq ~#q ~#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#sq ~ L�:�Wuq ~ O   q ~t bayw  Nsq ~ '�osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~#"q ~#!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#(sq ~ LD�]uq ~ O   q ~	q ~	w  Lsq ~ '&x�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt arlington_txt arlington_tx:cxq ~#/q ~#.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#8sq ~ L�Q��uq ~ O   q ~�q ~w  sq ~ 'FC�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(xq ~#?q ~#>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#Esq ~ Lf�4Fuq ~ O   q ~3t nhw  sq ~ '�,�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~#Mq ~#Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#Ssq ~ L��K5uq ~ O   q ~ Qq ~ Rq ~ Sq ~ gw  sq ~ '��fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Txq ~#Zq ~#Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#`sq ~ LJC@�uq ~ O   q ~ Qq ~ �q ~ q ~=w  	�sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t pearl_rivert pearl_river:rxq ~#gq ~#fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#psq ~ L���uq ~ O   q ~ Qt pearlw  sq ~ 'k��"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_rochelle_nyt new_rochelle_ny:cxq ~#xq ~#wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L0o�quq ~ O   q ~�t rochelleq ~�q ~�w  {sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L�!9uq ~ O   q ~�q ~Uw  �sq ~ ':�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~6t 	oakland:nxq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L�p*�uq ~ O   q ~6w  �sq ~ '�#��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L��)uq ~ O   q ~ �q ~q ~ �w  osq ~ '��#rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L'�uq ~ O   q ~Nq ~w  3sq ~ '%��-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L)��uq ~ O   q ~�w  sq ~ '�xj�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t wabash_rivert wabash_river:rxq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ LO*I�uq ~ O   q ~ Qt wabashq ~ �w  lsq ~ '-3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t kenner:nxq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L�Y{uq ~ O   q ~�w  sq ~ 'a#��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\xq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~#�sq ~ L2���uq ~ O   q ~ Rq ~ Sq ~�q ~4w  qsq ~ '>��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t silver_springt silver_spring:nxq ~#�q ~#�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$sq ~ LG_��uq ~ O   t silvert springw   �sq ~ '��+Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt whittier_cat whittier_ca:cxq ~$q ~$
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$sq ~ L~`>�uq ~ O   q ~�q ~"w  �sq ~ '
G��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~$q ~$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$!sq ~ L՛�(uq ~ O   q ~"w  �sq ~ 'G��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(xq ~$(q ~$'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$.sq ~ L�oӜuq ~ O   q ~ Qq ~ �q ~3q ~	bw  �sq ~ '��DJsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t cumberland_rivert cumberland_river:rxq ~$5q ~$4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$>sq ~ L��<uq ~ O   q ~ Qt 
cumberlandq ~ �w  *sq ~ 'e�V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~$Fq ~$Esq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~$Lsq ~ L��tjuq ~ O   t borderw   (sq ~ '� s�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~$Tq ~$Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$Zsq ~ L�5�Kuq ~ O   q ~�q ~
�q ~�w  	~sq ~ '�1�Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~$aq ~$`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$gsq ~ L�� �uq ~ O   q ~ Qq ~ �q ~�w  `sq ~ '���tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_mateo_cat san_mateo_ca:cxq ~$nq ~$msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$wsq ~ L�2&Luq ~ O   q ~ �t mateoq ~"w  }sq ~ '�'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cleveland_oht cleveland_oh:cxq ~$q ~$~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L��)uq ~ O   t 	clevelandq ~�w  �sq ~ '�'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt long_beach_cat long_beach_ca:cxq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L�nGuq ~ O   t longq ~	bw  Rsq ~ '�%M�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	orange_cat orange_ca:cxq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L��&luq ~ O   q ~hw  �sq ~ '0>�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Cxq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L�IDuq ~ O   q ~ Nw  %sq ~ 'p�tXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~<t portsmouth:nxq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L.� 3uq ~ O   q ~<w  �sq ~ '��3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt berkeley_cat berkeley_ca:cxq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L�
!uq ~ O   q ~�q ~"w  �sq ~ '��@�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L)��Zuq ~ O   q ~�w  Csq ~ 'aqCSsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~$�sq ~ L��uq ~ O   q ~�q ~	bq ~"w  �sq ~ ':�l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t equalst equals:<e,<e,t>>xq ~$�q ~$�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~% sq ~ Ld��Uuq ~ O   t 	excludingw   Gsq ~ '���5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt flint_mit 
flint_mi:cxq ~%q ~%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%sq ~ L~uq ~ O   q ~ Qq ~ �t flintw  sq ~ '�;��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#xq ~%q ~%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%sq ~ L�`��uq ~ O   q ~�q ~.w  )sq ~ '��9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~%&q ~%%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%,sq ~ LY4c�uq ~ O   q ~Cq ~�w  �sq ~ '��|8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
tuscaloosat tuscaloosa:nxq ~%3q ~%2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%<sq ~ L?j2�uq ~ O   q ~%5w  :sq ~ '�'usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~%Cq ~%Bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%Isq ~ L�~�'uq ~ O   q ~q ~"w  ysq ~ '�C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	boston_mat boston_ma:cxq ~%Pq ~%Osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%Ysq ~ L�Guq ~ O   t bostonq ~�w  �sq ~ 'h��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~cxq ~%aq ~%`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%gsq ~ L�5?8uq ~ O   q ~|q ~"w  	Asq ~ 'Yq�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t louisiana:sxq ~%nq ~%msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%vsq ~ L[ �uq ~ O   q ~ Rq ~ Sq ~�w  �sq ~ '�eY�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~%}q ~%|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ Lm�h�uq ~ O   q ~�q ~�q ~�w  �sq ~ '�ܪsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
 xq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ LV���uq ~ O   q ~
q ~
q ~w  sq ~ '�U�yq ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~%�q ~%�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~%�sq ~ LK�iuq ~ O   t 	traversesw  
sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt tuscaloosa_alt tuscaloosa_al:cxq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ Lv��uq ~ O   q ~%5q ~Iw  	hsq ~ '_�~dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt garden_grove_cat garden_grove_ca:cxq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ LUM	�uq ~ O   q ~q ~q ~ �w  sq ~ '6$rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ LS6^uq ~ O   q ~�q ~"w  �sq ~ '!/�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ L��r�uq ~ O   q ~q ~#q ~�w  sq ~ 'ߛssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bxq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ L�"�uq ~ O   q ~ Qq ~ �q ~Mw  (sq ~ '1+�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ L���uq ~ O   q ~Dq ~�w  	sq ~ '��9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~%�q ~%�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~%�sq ~ L�Nmuq ~ O   q ~�w  sq ~ 'm��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt waterford_mit waterford_mi:cxq ~&q ~&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&sq ~ LuImjuq ~ O   t 	waterfordq ~Tw  #sq ~ 'w\bxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~)t milwaukee:nxq ~&q ~&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&sq ~ L�>uq ~ O   q ~)w  �sq ~ '0��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~&#q ~&"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&)sq ~ L����uq ~ O   q ~ Qq ~�q ~ �w  �sq ~ '.H�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~&0q ~&/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&6sq ~ L��Tuq ~ O   q ~ Qq ~ �q ~�w  �sq ~ 'ʃ�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%oxq ~&=q ~&<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&Csq ~ L~l�uq ~ O   q ~�w  �sq ~ '�ػAsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~&Jq ~&Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&Psq ~ Lׯ��uq ~ O   q ~Dq ~�w  �sq ~ 'u��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt baltimore_mdt baltimore_md:cxq ~&Wq ~&Vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&`sq ~ L6�>�uq ~ O   q ~�t mdw  �sq ~ '��+�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt oklahoma_city_okt oklahoma_city_ok:cxq ~&hq ~&gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&qsq ~ L��uq ~ O   q ~�q ~ �q ~�w  Ksq ~ '�&��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t dundalkt 	dundalk:nxq ~&xq ~&wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ Lw�.wuq ~ O   q ~&zw  3sq ~ '��xPsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt waco_txt 	waco_tx:cxq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ LL�uq ~ O   t wacoq ~ �w  �sq ~ 'Іf�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
lincoln_net lincoln_ne:cxq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ L��uq ~ O   q ~ Qq ~ �t lincolnw  �sq ~ 'a�j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ixq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ Ly�&�uq ~ O   q ~�q ~tq ~�w  sq ~ '�Y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Wt 
amarillo:nxq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ L�W%uq ~ O   q ~Ww  Gsq ~ '%�Xcq ~�sq ~ sq ~ sq ~ J   w   q ~Aq ~�q ~�xq ~&�q ~&�sq ~ @q ~�sq ~ G���    sq ~ sq ~ J   w   q ~ �q ~q ~xq ~&�sq ~ L��$guq ~ O   t longerw  
?sq ~ 'vg~sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cherry_hill_njt cherry_hill_nj:cxq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ L�&�8uq ~ O   t cherryq ~�q ~�q ~Fw  9sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt somerville_mat somerville_ma:cxq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ L�Ruq ~ O   q ~!)w  �sq ~ '���csq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	joliet_ilt joliet_il:cxq ~&�q ~&�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~&�sq ~ LU���uq ~ O   t jolietq ~Uw  :sq ~ 'Nj��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	durham_nct durham_nc:cxq ~'q ~'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'sq ~ L�J�1uq ~ O   t durhamw  �sq ~ '��*_sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~'q ~'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'sq ~ L�ɫuq ~ O   q ~q ~.w  sq ~ '�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~'!q ~' sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~''sq ~ Ly���uq ~ O   q ~q ~�w  Nsq ~ '?Ce+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t ontariot 	ontario:lxq ~'.q ~'-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'7sq ~ L�8�=uq ~ O   q ~q ~'0w  Psq ~ 'dx�3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
memphis_tnt memphis_tn:cxq ~'>q ~'=sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'Gsq ~ LD͡uq ~ O   q ~ Qq ~ �t memphisw  �sq ~ '�fF�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
hammond_int hammond_in:cxq ~'Oq ~'Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'Xsq ~ Lr��uq ~ O   t hammondq ~iw  �sq ~ 'hחsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
lubbock_txt lubbock_tx:cxq ~'`q ~'_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'isq ~ L*���uq ~ O   q ~ Qq ~ �t lubbockw  	sq ~ '�I��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt erie_pat 	erie_pa:cxq ~'qq ~'psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'zsq ~ L /��uq ~ O   t eriew  Ysq ~ 'y+v3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t canadian_rivert canadian_river:rxq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ Lf��uq ~ O   t canadianq ~ �w  sq ~ 'x.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t greenville:nxq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ L�Nmuq ~ O   q ~�w  sq ~ '�&H[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ L�j{kuq ~ O   q ~wq ~�w  Gsq ~ '�b��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ L�0�uq ~ O   q ~!)q ~�w  gsq ~ '��3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt newport_news_vat newport_news_va:cxq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ LS9`�uq ~ O   q ~3t newsw  	sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt mountain_view_cat mountain_view_ca:cxq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ L4@~uq ~ O   q ~�q ~�q ~"w  �sq ~ '/�,`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ L���tuq ~ O   q ~�q ~�w  Esq ~ '��psq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
meriden_ctt meriden_ct:cxq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~'�sq ~ L8�huq ~ O   t meridenw  	]sq ~ '�>R!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~:xq ~'�q ~'�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ LIw@uq ~ O   q ~Ew  �sq ~ 'Mrsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~(q ~(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ L
H�uq ~ O   q ~ Qq ~ �q ~Cw  �sq ~ '��5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~(q ~(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ L���Juq ~ O   q ~Xq ~ �w  �sq ~ '$���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
yonkers_nyt yonkers_ny:cxq ~("q ~(!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(+sq ~ Lд��uq ~ O   q ~ Qq ~ �t yonkersw  �sq ~ '>|Jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~(3q ~(2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(9sq ~ LPw��uq ~ O   q ~ Qq ~ �q ~q ~w  5sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~(@q ~(?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(Fsq ~ LL'uq ~ O   q ~q ~Iw   �sq ~ 'S��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t oklahoma_cityt oklahoma_city:nxq ~(Mq ~(Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(Vsq ~ L��:uq ~ O   q ~�q ~ �w  �sq ~ '+w+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ gt 
michigan:lxq ~(]q ~(\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(esq ~ L�H�}uq ~ O   q ~q ~ gw  +sq ~ '�E1Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~(lq ~(ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(rsq ~ L�|��uq ~ O   q ~ Qq ~ �q ~&w  �sq ~ ';��,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~cxq ~(yq ~(xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(sq ~ L�j,�uq ~ O   q ~ Qq ~ �q ~nq ~w   �sq ~ 'P��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	escondidot escondido:nxq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ La��"uq ~ O   q ~(�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ L66
�uq ~ O   q ~�t njw  wsq ~ '[us;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ L$�<uq ~ O   q ~�q ~Mw  [sq ~ '�vbsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ L�{RQuq ~ O   q ~�q ~w  xsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'?xq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ L�Q��uq ~ O   q ~'Jq ~5w  �sq ~ '6�V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt south_bend_int south_bend_in:cxq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ LE�%Fuq ~ O   q ~ Qq ~ �q ~
�t bendw  �sq ~ '�#�q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~(�q ~(�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~(�sq ~ L���uq ~ O   q ~�w  

sq ~ '��dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt jersey_city_njt jersey_city_nj:cxq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ L"���uq ~ O   q ~Fq ~ �q ~�q ~Fw  sq ~ 'w�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	denver_cot denver_co:cxq ~(�q ~(�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~(�sq ~ L7Гuq ~ O   t denverq ~#w  sq ~ '��9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lower_merion_pat lower_merion_pa:cxq ~)q ~)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)sq ~ LN �uq ~ O   t lowert merionq ~�w  lsq ~ ';��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~)q ~)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)sq ~ L�:�#uq ~ O   q ~+q ~�w  zsq ~ 'g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	hxq ~)&q ~)%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~),sq ~ L�-:uq ~ O   q ~�q ~	sq ~Uw  �sq ~ '6�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
dubuque_iat dubuque_ia:cxq ~)3q ~)2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)<sq ~ Lox�uq ~ O   t dubuqueq ~ w  Csq ~ 'J�~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~)Dq ~)Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)Jsq ~ L;p�uq ~ O   q ~ Qq ~ �q ~<w  sq ~ '00q ~�sq ~ sq ~ sq ~ J   w   q ~Zxq ~)Pq ~)Osq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)Tsq ~ L9W�uq ~ O   t countryw  
2sq ~ 'j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~)\q ~)[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)bsq ~ L=b�uq ~ O   q ~�w  jsq ~ '�?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~)iq ~)hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)osq ~ L#���uq ~ O   q ~�w  �sq ~ '�?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t little_missouri_rivert little_missouri_river:rxq ~)vq ~)usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)sq ~ Lɏ:uq ~ O   q ~ Qq ~�q ~�w  \sq ~ '��׭sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L�,S�uq ~ O   q ~�w  �sq ~ ' �{{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ LIj��uq ~ O   q ~!)q ~�w  �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t brownsville:nxq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L�sóuq ~ O   q ~�w  sq ~ 'r�<-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L���uq ~ O   q ~�q ~�q ~Fw  ksq ~ 'ꪓ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt san_antonio_txt san_antonio_tx:cxq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L;�uq ~ O   q ~ �t antoniow  =sq ~ '�՝Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L�{�uq ~ O   q ~�w  �sq ~ 'L�"Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ LA�Zuq ~ O   q ~Mw  �sq ~ '��I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L���uq ~ O   q ~ Qq ~ Rq ~ Sq ~Uq ~�w  �sq ~ ' ��}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt honolulu_hit honolulu_hi:cxq ~)�q ~)�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~)�sq ~ L{�+)uq ~ O   q ~ q ~w  8sq ~ '�װ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	redford:nxq ~*q ~*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*sq ~ L@�
uq ~ O   q ~�w  .sq ~ 'ѬNXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t cheektowagat cheektowaga:nxq ~*q ~*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*sq ~ L5�C#uq ~ O   q ~*w  �sq ~ '� ]zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt boise_idt 
boise_id:cxq ~*#q ~*"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*,sq ~ L�Luq ~ O   q ~�w   �sq ~ '�k�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%�xq ~*3q ~*2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*9sq ~ LuS�8uq ~ O   q ~ Qq ~ �q ~q ~w   �sq ~ '�MJ3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t 	montana:sxq ~*@q ~*?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*Hsq ~ L�uq ~ O   q ~�q ~ Rw   �sq ~ '�^�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt ann_arbor_mit ann_arbor_mi:cxq ~*Oq ~*Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*Xsq ~ LM���uq ~ O   t annt arborq ~ gw  	_sq ~ 'K|)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~*aq ~*`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*gsq ~ LOn_iuq ~ O   q ~ fq ~�q ~Tw  �sq ~ 'd��5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	irvine_cat irvine_ca:cxq ~*nq ~*msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*wsq ~ L[��uq ~ O   t irvineq ~"w  �sq ~ 'PLزsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~cxq ~*q ~*~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ L�|+uq ~ O   q ~nq ~q ~"w  �sq ~ 'H���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ L�Kuq ~ O   q ~Dq ~Ew  �sq ~ '��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
alhambra:nxq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ Ldt�&uq ~ O   q ~�w  �sq ~ '�'�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_alverstonet mount_alverstone:mxq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ Lf�z�uq ~ O   q ~ zt 
alverstonew  Ksq ~ 'XH��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ L��Vuq ~ O   q ~ �w  sq ~ ' L�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~*�sq ~ L �]uq ~ O   t youw  	�sq ~ '�7�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ L�0��uq ~ O   q ~&�w  �sq ~ '1>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ L
���uq ~ O   q ~ Qq ~ �q ~Dw  	�sq ~ '	�B+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~*�sq ~ Lm���uq ~ O   q ~�q ~ gw  �sq ~ ' �sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~*�q ~*�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~*�sq ~ L ��uq ~ O   q ~w   sq ~ ':�$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~+q ~+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+	sq ~ L݇�uq ~ O   q ~�q ~ �w  �sq ~ 'Ҡu5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
burbank_cat burbank_ca:cxq ~+q ~+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+sq ~ L����uq ~ O   q ~ �q ~"w  �sq ~ '���q ~�sq ~ sq ~ sq ~ J   w   q ~Hq ~Hxq ~+q ~+sq ~ @q ~�sq ~ Go��    sq ~ sq ~ J   w   q ~q ~xq ~+#sq ~ L�p
uq ~ O   q ~Sw  	�sq ~ '=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~+*q ~+)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+0sq ~ L9�"cuq ~ O   q ~ Rq ~ Sq ~Uw  |sq ~ '��tMsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<xq ~+7q ~+6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+=sq ~ L���uq ~ O   q ~ Qq ~ �q ~Gw  esq ~ 'qE<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
louisvillet louisville:nxq ~+Dq ~+Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+Msq ~ LO�-uq ~ O   q ~+Fw  sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t alaskat alaska:nxq ~+Tq ~+Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+]sq ~ L����uq ~ O   q ~+Vw  �sq ~ 'WE��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~+dq ~+csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+jsq ~ L���uq ~ O   q ~ Qq ~ �q ~q ~q ~ �w  �sq ~ '7�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
medford_mat medford_ma:cxq ~+qq ~+psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+zsq ~ LDJ]+uq ~ O   q ~ Qq ~ �t medfordw  �sq ~ 'w��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	pomona_cat pomona_ca:cxq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ L�X	juq ~ O   t pomonaq ~ �w  	�sq ~ '��Y�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ L���uq ~ O   q ~�q ~Ew   tsq ~ '�YZq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~+�sq ~ L�X�uq ~ O   q ~"w  
1sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ LH���uq ~ O   q ~'�q ~�w  �sq ~ '~�> sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*xq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ L��<tuq ~ O   q ~ q ~5w  �sq ~ '���|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t connecticut_rivert connecticut_river:rxq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ Lg��uq ~ O   q ~ Qq ~�w  ;sq ~ 'ĩ�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~	�t new_mexico:nxq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ L��2�uq ~ O   q ~�q ~�w  �sq ~ 'ꈐsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt scranton_pat scranton_pa:cxq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ L�C3buq ~ O   t scrantonw  fsq ~ '�cV\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Cxq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~+�sq ~ L����uq ~ O   q ~ Nq ~�w  Hsq ~ '��u�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~+�q ~+�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,sq ~ L쮫�uq ~ O   q ~ �q ~Nq ~"w  Isq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
vallejo_cat vallejo_ca:cxq ~,q ~,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,sq ~ L_�uq ~ O   q ~ Qq ~ �t vallejow  �sq ~ '01Q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~,q ~,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,#sq ~ Lc.s�uq ~ O   q ~ Qq ~ Rq ~ Sq ~q ~ w  sq ~ '�msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(#xq ~,*q ~,)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,0sq ~ L��c uq ~ O   q ~(.q ~�q ~�w  �sq ~ '��(Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~,7q ~,6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,=sq ~ LM�5�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��l{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
new_york:nxq ~,Dq ~,Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,Lsq ~ L l>uq ~ O   q ~�q ~�w  6sq ~ '��z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~,Sq ~,Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,Ysq ~ L��7�uq ~ O   q ~	�w  �sq ~ '�7�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~,`q ~,_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,fsq ~ L Ӓ�uq ~ O   q ~�q ~	�w  �sq ~ '�M��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~,mq ~,lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,ssq ~ L
��=uq ~ O   q ~&�w  ^sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
ontario_cat ontario_ca:cxq ~,zq ~,ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ L�t�uq ~ O   q ~'0q ~ �w  sq ~ '��g�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt escondido_cat escondido_ca:cxq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ L�)4uq ~ O   q ~(�q ~"w  sq ~ '{���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ L���\uq ~ O   q ~	�q ~�w   �sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ LFɐxuq ~ O   q ~&�t new  sq ~ 'R�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt glendale_azt glendale_az:cxq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ Lۈ��uq ~ O   q ~ Qq ~ �t glendalew  �sq ~ '�t��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t canton:nxq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ L�zo�uq ~ O   q ~�w  Osq ~ 'w��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~,�sq ~ L 7�uq ~ O   q ~w   Msq ~ 'rJ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ L<e_�uq ~ O   q ~ Qq ~ �q ~Hw  �sq ~ 'U�L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~,�sq ~ L'B`�uq ~ O   q ~�q ~�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~,�q ~,�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-sq ~ L.��uq ~ O   q ~ Qq ~ �q ~�q ~�w  sq ~ '�|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~-	q ~-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-sq ~ LC�8uq ~ O   q ~ Qq ~ �q ~q ~ �w  6sq ~ 'n��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~-q ~-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~-sq ~ L 3;�uq ~ O   q ~w   )sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~-#q ~-"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-)sq ~ LΉ�
uq ~ O   q ~qq ~ �w  sq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~nxq ~-0q ~-/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-6sq ~ L�"�uq ~ O   q ~yq ~ �w  lsq ~ '�S �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt alexandria_vat alexandria_va:cxq ~-=q ~-<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-Fsq ~ L�p�uq ~ O   q ~ Qq ~ �q ~�w  $sq ~ 'Z�m�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt woodbridge_njt woodbridge_nj:cxq ~-Mq ~-Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-Vsq ~ L��4Duq ~ O   t 
woodbridgeq ~�q ~Fw   �sq ~ 'p3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~-^q ~-]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-dsq ~ L�iUuq ~ O   q ~ Qq ~ �q ~&�w  %sq ~ '	:�ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~-kq ~-jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-qsq ~ Lrduq ~ O   q ~&q ~ gw  �sq ~ 'Ӊ&8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t greensboro:nxq ~-xq ~-wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L���Xuq ~ O   q ~�w  isq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	oxnard_cat oxnard_ca:cxq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L�p�2uq ~ O   q ~ Qq ~ �t oxnardw  	�sq ~ '��&sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~-�sq ~ L�C�uq ~ O   t tellt mew   sq ~ '<��q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~-�q ~-�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~-�sq ~ L  cuq ~ O   q ~w  	�sq ~ '  ��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~-�sq ~ L  �uq ~ O   t kmw  	�sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~+Vt alaska:sxq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L:�ًuq ~ O   q ~ Rq ~ Sq ~+Vw  
sq ~ '��Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L�d�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��^]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	pueblo_cot pueblo_co:cxq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L��[	uq ~ O   q ~ Qq ~ �t pueblow  /sq ~ '���[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L�{��uq ~ O   q ~Dq ~	�w  �sq ~ 'م�@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt evansville_int evansville_in:cxq ~-�q ~-�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-�sq ~ L/\��uq ~ O   t 
evansvilleq ~iw  Usq ~ 'ɍ_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
costa_mesat costa_mesa:nxq ~.q ~.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.sq ~ L�uuq ~ O   q ~�q ~�w  �sq ~ '�"8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Xt 
columbia:nxq ~.q ~.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.sq ~ L��6 uq ~ O   q ~Xw  �sq ~ '��I�q ~�sq ~ sq ~ sq ~ J   w   q ~xq ~.#q ~."sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~.'sq ~ L 2�*uq ~ O   t livew  	�sq ~ '��6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	detroit:nxq ~./q ~..sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.7sq ~ L\���uq ~ O   q ~�w  	.sq ~ '��ğsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%Qxq ~.>q ~.=sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.Dsq ~ L��&uq ~ O   q ~%\w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt syracuse_nyt syracuse_ny:cxq ~.Kq ~.Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.Tsq ~ L?�}uq ~ O   q ~ Qq ~ �t syracusew  �sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~.\q ~.[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.bsq ~ L�Wz�uq ~ O   q ~�q ~`w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%oxq ~.iq ~.hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.osq ~ LU�&�uq ~ O   q ~�q ~ Rw  �sq ~ '1�!gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_hubbardt mount_hubbard:mxq ~.vq ~.usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.sq ~ Lduq ~ O   q ~ zt hubbardw  �sq ~ '�X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt bethlehem_pat bethlehem_pa:cxq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ LP�
quq ~ O   t 	bethlehemq ~�w  �sq ~ '�W��q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ �M�t <l,t>q ~�q ~ �q ~t 
lake:<l,t>xq ~.�q ~.�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~.�sq ~ L�uq ~ O   t lakesw  	�sq ~ '�X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*$xq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ L�}�uq ~ O   q ~ Qq ~ �q ~�w  	vsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ LսU^uq ~ O   q ~�q ~�q ~w  *sq ~ ')��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt east_orange_njt east_orange_nj:cxq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ Li�z�uq ~ O   q ~gq ~hq ~(�w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ L��]uq ~ O   q ~�q ~	bq ~ �w   �sq ~ '���rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ L,khuq ~ O   q ~ Rq ~ Sq ~�w  	2sq ~ '�0Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt springfield_mot springfield_mo:cxq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~.�sq ~ L��uq ~ O   q ~Fq ~�w  sq ~ 'CR�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~.�q ~.�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/sq ~ L��uq ~ O   q ~�w  �sq ~ 'X���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
clinton_mit clinton_mi:cxq ~/q ~/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/sq ~ L6���uq ~ O   t clintonq ~Tw  �sq ~ 'I�!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Axq ~/q ~/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/sq ~ LE���uq ~ O   q ~Lq ~Iw  �sq ~ '1�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~/&q ~/%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/,sq ~ L�@��uq ~ O   q ~5w  dsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t south_carolinat south_carolina:sxq ~/3q ~/2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/<sq ~ L�F�uq ~ O   q ~ Rq ~ Sq ~
�q ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~/Cq ~/Bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/Isq ~ L[��uq ~ O   q ~7t hiw  �sq ~ 'ZZ.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~/Qq ~/Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/Wsq ~ LFfR�uq ~ O   q ~ Qq ~ �q ~�w  sq ~ '�;D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~/^q ~/]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/dsq ~ LY�!+uq ~ O   q ~�w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~/kq ~/jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/qsq ~ L~d$�uq ~ O   q ~)q ~)w  osq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt inglewood_cat inglewood_ca:cxq ~/xq ~/wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ L�}��uq ~ O   t 	inglewoodq ~"w  :sq ~ 't�k�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+xq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ L��(�uq ~ O   q ~6q ~"w  	asq ~ '�Wcsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ L�u�uq ~ O   q ~ Qq ~ Rq ~ Sq ~w  �sq ~ '	 �dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#xq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ LF/�uq ~ O   q ~�q ~.q ~�w  �sq ~ '�$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
norfolk_vat norfolk_va:cxq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ L�V�uq ~ O   q ~ Qq ~ �t norfolkw  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ L�9�uq ~ O   q ~"	q ~(�w  =sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t westminster:nxq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ L���uq ~ O   q ~w  Ksq ~ '?�:vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t republican_rivert republican_river:rxq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ LTRuq ~ O   q ~ Qt 
republicanq ~ �w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~{xq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/�sq ~ Lp|�uq ~ O   q ~�q ~�w  sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~/�q ~/�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0sq ~ L�L�Quq ~ O   q ~
Yq ~ �w  xsq ~ '�Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt chesapeake_vat chesapeake_va:cxq ~0q ~0sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0sq ~ L($��uq ~ O   t 
chesapeakeq ~ w  �sq ~ '�3�jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&Xxq ~0q ~0sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0sq ~ LF>�ouq ~ O   q ~�q ~�w  Ssq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~0&q ~0%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0,sq ~ L�mR8uq ~ O   q ~�q ~Eq ~�q ~�w  =sq ~ 'a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt evanston_ilt evanston_il:cxq ~03q ~02sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0<sq ~ L��Buq ~ O   q ~ Qq ~ �t evanstonw   ksq ~ '|z�Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
roanoke_vat roanoke_va:cxq ~0Dq ~0Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0Msq ~ LQz��uq ~ O   q ~<w  �sq ~ '�7(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt new_york_nyt new_york_ny:cxq ~0Tq ~0Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0]sq ~ L�~��uq ~ O   q ~ Qq ~ �q ~ Sq ~�q ~�w  ?sq ~ '�HH�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~0dq ~0csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0jsq ~ Lz�L�uq ~ O   q ~
�q ~
�w  }sq ~ '�O�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	6xq ~0qq ~0psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0wsq ~ L��xuq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  3sq ~ '�]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~0~q ~0}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ LR���uq ~ O   q ~�q ~�q ~Tw  �sq ~ ' �9�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~0�sq ~ L ���uq ~ O   q ~<w  
%sq ~ ' 8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~0�sq ~ L ��uq ~ O   q ~ Qw   sq ~ 'vU9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~ t 
virginia:sxq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ L\�Mcuq ~ O   q ~ w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Yxq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ L��:!uq ~ O   q ~ fq ~Tw  �sq ~ 'E�K�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ Lb�B�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ 'M˗�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt nashville_tnt nashville_tn:cxq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ L�.�uq ~ O   t 	nashvillet tnw  4sq ~ '? ԛsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~/5t south_carolina:nxq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ Lʸ�>uq ~ O   q ~
�q ~�w  �sq ~ '  q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~0�sq ~ L  �uq ~ O   t 50w  
sq ~ 'Qʣ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_castlet mount_castle:mxq ~0�q ~0�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~0�sq ~ Ln���uq ~ O   q ~ zt castlew  �sq ~ '3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt louisville_kyt louisville_ky:cxq ~1q ~1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1sq ~ L����uq ~ O   q ~+Fq ~Mw  �sq ~ 'J;,q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~1q ~1sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~1sq ~ L�Z�2uq ~ O   t flowingw  
8sq ~ '�Ouq ~�sq ~ sq ~ sq ~ J   w   q ~xq ~1q ~1sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~1"sq ~ L�v�uq ~ O   t therew  
sq ~ 'ǕW�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~1*q ~1)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~10sq ~ L�Y�duq ~ O   q ~ Qq ~ �q ~�w  	Dsq ~ '�.;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt winston-salem_nct winston-salem_nc:cxq ~17q ~16sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1@sq ~ L�۾`uq ~ O   t winston-salemq ~_w  �sq ~ '5�~+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t huront huron:lxq ~1Hq ~1Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1Qsq ~ L�uq ~ O   q ~q ~1Jw  sq ~ '8S�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*Axq ~1Xq ~1Wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1^sq ~ L����uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w   �sq ~ '8UU[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_biancat mount_bianca:mxq ~1eq ~1dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1nsq ~ Lm���uq ~ O   q ~ zt biancaw  �sq ~ '�Q��q ~�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~t 0t 0:ixq ~1uq ~1tsq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1|q ~�w   Lsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ >t maine:nxq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L-�
uq ~ O   q ~ >w  �sq ~ '��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L�kg�uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  4sq ~ '�'	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t ouachita_rivert ouachita_river:rxq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L�$��uq ~ O   t ouachitaq ~ �w  �sq ~ '�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t topekat topeka:nxq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L�B�Duq ~ O   q ~1�w  0sq ~ '8��q ~�sq ~ sq ~ sq ~ J   w   q ~:xq ~1�q ~1�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~1�sq ~ L���@uq ~ O   q ~!�w  
sq ~ '!	��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~)t denver:nxq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L�g��uq ~ O   q ~)w  �sq ~ '�z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
el_paso_txt el_paso_tx:cxq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L 5�&uq ~ O   q ~ �t pasow  �sq ~ '��a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ LO�-uq ~ O   q ~+Fw  sq ~ '�ʡ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~1�q ~1�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~1�sq ~ L�f�uq ~ O   q ~ Qq ~ �q ~	q ~	w  sq ~ 'y�}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Txq ~2q ~2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2sq ~ L�m�zuq ~ O   q ~ q ~=w  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~2q ~2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2sq ~ L ?��uq ~ O   q ~ Qq ~ Rq ~ Sq ~�q ~�w  'sq ~ 'JS6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~&t odessa:nxq ~2q ~2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2$sq ~ L��uq ~ O   q ~&w  �sq ~ 'YX# sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_la_platat mount_la_plata:mxq ~2+q ~2*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~24sq ~ LPt��uq ~ O   q ~ zq ~"�t plataw  jsq ~ 'P�%5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~2<q ~2;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2Bsq ~ L�+T=uq ~ O   q ~�q ~"w  �sq ~ '�@v'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_fairweathert mount_fairweather:mxq ~2Iq ~2Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2Rsq ~ L��7uq ~ O   q ~ zt fairweatherw  �sq ~ '�*�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#yxq ~2Zq ~2Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2`sq ~ L[��\uq ~ O   q ~ Qq ~ �q ~�q ~#�w  osq ~ '�a&sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~2gq ~2fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2msq ~ L�zo�uq ~ O   q ~�w  �sq ~ '�.�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~2tq ~2ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2zsq ~ L�h�~uq ~ O   q ~q ~(�w  /sq ~ '�]bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~dxq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ LM�WEuq ~ O   q ~ Qq ~ �q ~oq ~pw  �sq ~ '  �Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~2�sq ~ L  uq ~ O   q ~ Sw   +sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t el_cajont 
el_cajon:nxq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ L�V�uq ~ O   q ~ �q ~ �w  Asq ~ '�+�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt pawtucket_rit pawtucket_ri:cxq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ L��uq ~ O   q ~ Qq ~ �t 	pawtucketw  �sq ~ '�<�1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ LEE�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��٤sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~2�sq ~ L��aeuq ~ O   q ~t metersw   sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
waltham_mat waltham_ma:cxq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ L�P_<uq ~ O   t walthamq ~�w  �sq ~ '�p�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt levittown_nyt levittown_ny:cxq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ L����uq ~ O   t 	levittownw  Ssq ~ 'o�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~2�q ~2�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~2�sq ~ L��uq ~ O   q ~Hq ~Mw  �sq ~ '��$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0Exq ~3q ~3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3sq ~ L]�WCuq ~ O   q ~ Qq ~ �q ~<w  hsq ~ 'ZC�%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt lawrence_mat lawrence_ma:cxq ~3q ~3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3sq ~ L
�uq ~ O   q ~~q ~�w  	�sq ~ '/�o�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~3#q ~3"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3)sq ~ L�4Huuq ~ O   q ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~30q ~3/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~36sq ~ L���%uq ~ O   q ~�q ~�w  �sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~3=q ~3<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3Csq ~ L|�<huq ~ O   q ~ Qq ~ �q ~
w  �sq ~ '��+<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/�xq ~3Jq ~3Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3Psq ~ L�Euq ~ O   q ~ Qq ~/�w  Ysq ~ '�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~3Wq ~3Vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3]sq ~ L,ףyuq ~ O   q ~ Qq ~ �q ~Nw  usq ~ 'CZ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~3dq ~3csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3jsq ~ L�J(|uq ~ O   q ~Dq ~iw  esq ~ '���xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t rockfordt 
rockford:nxq ~3qq ~3psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3zsq ~ L�Q�uq ~ O   q ~3sw   �sq ~ '�4�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~vxq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ L�<�uq ~ O   q ~�q ~*w   �sq ~ 'c$�%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ L+��+uq ~ O   q ~�q ~�w  (sq ~ '�Yڃsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ L���5uq ~ O   q ~ Qq ~ �q ~w  	 sq ~ 'ꃈ+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ Lc�\�uq ~ O   q ~�q ~�w  �sq ~ '�*�csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0�xq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ L�s�uq ~ O   q ~ Qq ~ Rq ~ Sq ~ w  	�sq ~ 'Uj�:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!uxq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ Ldo�uq ~ O   q ~ �q ~!�q ~ �w   �sq ~ '$�+�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ L��b�uq ~ O   q ~�q ~Iw  1sq ~ '��0�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~{xq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ Lj݌�uq ~ O   q ~ Qq ~ �q ~�w  [sq ~ '7o�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt buena_park_cat buena_park_ca:cxq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~3�sq ~ L���uq ~ O   t buenaq ~pq ~"w  7sq ~ '��=5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
trenton_njt trenton_nj:cxq ~3�q ~3�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4sq ~ L��X�uq ~ O   q ~�w  Vsq ~ '�^ktsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~4
q ~4	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4sq ~ Loe4�uq ~ O   q ~ q ~$q ~ �w  	Lsq ~ 'g�}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt 
mount_bonat mount_bona:mxq ~4q ~4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4 sq ~ L����uq ~ O   q ~ zt bonaw  Qsq ~ 'yl��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~4(q ~4'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4.sq ~ L�Ruq ~ O   q ~�q ~"�w  sq ~ '�\�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,{xq ~45q ~44sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4;sq ~ L�=Juq ~ O   q ~'0w  �sq ~ 'W�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ft 
stockton:nxq ~4Bq ~4Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4Jsq ~ Le�j�uq ~ O   q ~Fw  sq ~ '�$ōsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0Uxq ~4Qq ~4Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4Wsq ~ L l>uq ~ O   q ~�q ~�w  xsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~4^q ~4]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4dsq ~ L8��^uq ~ O   q ~�w  Ksq ~ '�y[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~wxq ~4kq ~4jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4qsq ~ L���uq ~ O   q ~�q ~q ~ w  2sq ~ '�N� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~4xq ~4wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4~sq ~ L�^uq ~ O   q ~ �q ~xw  	�sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(#xq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ L�
��uq ~ O   q ~(.q ~�w  bsq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt silver_spring_mdt silver_spring_md:cxq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ L��$uq ~ O   q ~$q ~$q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t redondo_beacht redondo_beach:nxq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ Lפ�uq ~ O   q ~	aq ~	bw  �sq ~ '�i8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ LĪ�uq ~ O   q ~ Qq ~ �q ~�w  +sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~dxq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ L��;uq ~ O   q ~oq ~pq ~�w  �sq ~ '϶\Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*xq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ L�Z�uq ~ O   q ~ q ~5q ~ �w  	jsq ~ '�{Q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ L��uq ~ O   q ~ Qq ~ �q ~)w  �sq ~ '�-8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~2�t 	waltham:nxq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ LB���uq ~ O   q ~2�w  ]sq ~ 'K��Zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#xq ~4�q ~4�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~4�sq ~ LY��vuq ~ O   q ~�q ~.q ~�w  	!sq ~ 'd��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4xq ~5q ~5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5sq ~ L��3uq ~ O   q ~?w  �sq ~ '��S�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t south_platte_rivert south_platte_river:rxq ~5q ~5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5sq ~ L<o�Huq ~ O   q ~ Qq ~
�t platteq ~ �w  �sq ~ '�s{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~pxq ~5 q ~5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5&sq ~ L[�'duq ~ O   q ~{q ~ �w  �sq ~ 'UAX�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~5-q ~5,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~53sq ~ L�?-�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ 'g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~5:q ~59sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~5@sq ~ L�+X�uq ~ O   t biggestw   sq ~ '�@Exsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~5Hq ~5Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5Nsq ~ L>6��uq ~ O   q ~q ~ �q ~�w  Esq ~ 'J«�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~5Uq ~5Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5[sq ~ L��uuq ~ O   q ~ q ~$w  �sq ~ '-��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t mississippi_rivert mississippi_river:rxq ~5bq ~5asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5ksq ~ Lߥ��uq ~ O   q ~�q ~ �w  �sq ~ '�}��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~5rq ~5qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5xsq ~ L�q�uq ~ O   q ~Hq ~Tw  :sq ~ '��$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	!xq ~5q ~5~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~5�sq ~ L��7,uq ~ O   t fewestw   %sq ~ 'w��q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~5�q ~5�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~5�sq ~ L 5��uq ~ O   t runsw  	�sq ~ '�"�'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ LpZuq ~ O   q ~ Qq ~ �q ~&�w  ^sq ~ '���ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ L	#|Luq ~ O   q ~ Qq ~ �q ~�w  sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~It 	alabama:sxq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ LW�ʁuq ~ O   q ~ Rq ~ Sq ~Iw  sq ~ 'FOsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,�xq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ L�P�Buq ~ O   q ~,�w  sq ~ '´sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Mxq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ L�|]5uq ~ O   q ~Xq ~�w  tsq ~ '�\Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	Vxq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ Lޯ�uq ~ O   q ~	aq ~	bq ~ �w  xsq ~ '
D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
penn_hillst penn_hills:nxq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ LD�]uq ~ O   q ~	q ~	w   �sq ~ 'i�ݩsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+xq ~5�q ~5�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~5�sq ~ L����uq ~ O   q ~ Qq ~ �q ~6w  	wsq ~ '<��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~6q ~6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6sq ~ La�?ruq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t west_hartfordt west_hartford:nxq ~6q ~6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6sq ~ L�pGuq ~ O   q ~q ~Cw  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt grand_rapids_mit grand_rapids_mi:cxq ~6"q ~6!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6+sq ~ L~KCKuq ~ O   q ~�q ~�w  sq ~ '�̸Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Wt oceanside:nxq ~62q ~61sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6:sq ~ L _�uq ~ O   q ~Ww  �sq ~ ' �?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~6Aq ~6@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6Gsq ~ L?���uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�QN{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
sioux_cityt sioux_city:nxq ~6Nq ~6Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6Wsq ~ L�gˏuq ~ O   q ~Uq ~ �w  sq ~ '�=Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~6^q ~6]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6dsq ~ L�{$uq ~ O   q ~ Qq ~ �q ~
�w   �sq ~ '��*sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~_xq ~6kq ~6jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6qsq ~ L,w�uq ~ O   q ~jw  	zsq ~ '�	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ixq ~6xq ~6wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6~sq ~ L܌+uq ~ O   q ~�q ~tw  �sq ~ '�rءsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
long_beacht long_beach:nxq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L�nGuq ~ O   q ~$�q ~	bw  Bsq ~ ' /�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~6�sq ~ L .��uq ~ O   q ~ �w  	�sq ~ 'd��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L����uq ~ O   q ~ Qq ~ �q ~ �w  �sq ~ '�>��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L �Vuq ~ O   q ~
�q ~(�q ~iw  sq ~ '�	Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L�jc_uq ~ O   q ~�w  sq ~ 'M�l8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~it 	indiana:nxq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ Ls��huq ~ O   q ~iw   �sq ~ '�/<5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt riverside_cat riverside_ca:cxq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L�E�uq ~ O   t 	riversideq ~"w  asq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L@_�uq ~ O   q ~ Qq ~ �q ~�q ~	bw   �sq ~ '�-8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6�sq ~ L�� uq ~ O   q ~�t nmw  �sq ~ '>�HUsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt washington_dct washington_dc:cxq ~6�q ~6�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7sq ~ L� s	uq ~ O   q ~�q ~Wq ~ Sq ~Xw  �sq ~ '�SUsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~7q ~7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7sq ~ L9^4�uq ~ O   q ~ Qq ~ �q ~ �w  �sq ~ 'R��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~7sq ~ LRNuq ~ O   t otherw  
5sq ~ '�Z�Fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~7%q ~7$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7+sq ~ L�Q�uq ~ O   q ~ Qq ~ �q ~�q ~�w  �sq ~ ')G8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~72q ~71sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~78sq ~ LL�suq ~ O   q ~�w  Zsq ~ '"=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fargo_ndt 
fargo_nd:cxq ~7?q ~7>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7Hsq ~ L1�fuq ~ O   t fargoq ~Uq ~
�w  �sq ~ 'H��_sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~7Pq ~7Osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7Vsq ~ LuSyuq ~ O   q ~[w  #sq ~ '��t�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
modesto_cat modesto_ca:cxq ~7]q ~7\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7fsq ~ L���uq ~ O   t modestoq ~ �w  Ksq ~ '��Ɵq ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~7mq ~7lsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~7qsq ~ L 2ƺuq ~ O   q ~$�w  	�sq ~ 'o�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	warren_mit warren_mi:cxq ~7xq ~7wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ LC�)uq ~ O   t warrenq ~Tw  �sq ~ '�p�Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~18xq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L~yuq ~ O   q ~ Qq ~ �q ~1Cw  	�sq ~ '�\�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t 
rock_rivert rock_river:rxq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L�k'uq ~ O   q ~�q ~ �w  Fsq ~ 'B���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L�*�juq ~ O   q ~wq ~�w  	sq ~ '���zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
decatur_ilt decatur_il:cxq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L[�Puq ~ O   t decaturw  	�sq ~ '0��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L�k4uq ~ O   q ~�q ~"w  �sq ~ '�
j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ LLt�uq ~ O   q ~ Qq ~ �q ~�q ~�w  �sq ~ '���[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%�xq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L��2�uq ~ O   q ~%5q ~Mw  �sq ~ '6P�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	Exq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ L|�Auq ~ O   q ~	Pq ~ �q ~�w   �sq ~ '�Ϭ{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~7�q ~7�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~7�sq ~ LQ7��uq ~ O   q ~�q ~�w  �sq ~ '�/��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~cxq ~8q ~8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8sq ~ L�(uq ~ O   q ~ Qq ~ �q ~|w  sq ~ '�4�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~8q ~8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8sq ~ L����uq ~ O   q ~Fq ~ �q ~(�w  fsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~8q ~8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8%sq ~ L��#uq ~ O   q ~ Qq ~ �q ~�w  sq ~ '�}vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt citrus_heights_cat citrus_heights_ca:cxq ~8,q ~8+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~85sq ~ L^��Juq ~ O   q ~�q ~�w  bsq ~ '�bFsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
midland_txt midland_tx:cxq ~8<q ~8;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8Esq ~ L�đuq ~ O   q ~�q ~w   �sq ~ '�<~sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t chattahoochee_rivert chattahoochee_river:rxq ~8Lq ~8Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8Usq ~ LE�7uq ~ O   q ~ Qt chattahoocheew  zsq ~ '�+	<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt ewa_hit ewa_hi:cxq ~8]q ~8\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8fsq ~ L9��uq ~ O   q ~ Qq ~ �t ewaw  sq ~ ' �(Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~~xq ~8nq ~8msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8tsq ~ L�Ԧuq ~ O   q ~�q ~�q ~ �w  �sq ~ 'j���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt manchester_nht manchester_nh:cxq ~8{q ~8zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ Ls)xuq ~ O   q ~ Qq ~ �t 
manchesterw  �sq ~ ' �gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_churchillt mount_churchill:mxq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L?��uq ~ O   q ~ zt 	churchillw  �sq ~ '�$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t pecos_rivert pecos_river:rxq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L�T��uq ~ O   t pecosq ~ �w  �sq ~ '@�G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt torrance_cat torrance_ca:cxq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L�ضuq ~ O   q ~!�w  <sq ~ ''��asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ LD��uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�Isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L�,ٸuq ~ O   q ~�w  �sq ~ '��`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L����uq ~ O   q ~ Qq ~ �q ~*w   �sq ~ '�X!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t chattanoogat chattanooga:nxq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L�X��uq ~ O   q ~8�w  Lsq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~et new_jersey:sxq ~8�q ~8�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~8�sq ~ L��B?uq ~ O   q ~�q ~Fq ~ Rw  �sq ~ 'fE�q ~�sq ~ sq ~ sq ~ J   w   q ~|xq ~9q ~9sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~9sq ~ L�l]!uq ~ O   t pointsw  	�sq ~ ')��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%	xq ~9q ~9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9sq ~ L�1�3uq ~ O   q ~%q ~Tw  �sq ~ '�vo[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~9q ~9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9"sq ~ L̕�Cuq ~ O   q ~�q ~�w  	"sq ~ '6��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~9)q ~9(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9/sq ~ L[4�uq ~ O   q ~�q ~5w  �sq ~ 'Yr	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0	xq ~96q ~95sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9<sq ~ LˆPSuq ~ O   q ~0q ~=w  Xsq ~ ''C�Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~9Cq ~9Bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9Isq ~ L�1�Kuq ~ O   q ~Fw  �sq ~ '�[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~9Pq ~9Osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9Vsq ~ L�|3�uq ~ O   q ~�w  Ysq ~ '�a��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t north_charlestont north_charleston:nxq ~9]q ~9\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9fsq ~ L#�Juq ~ O   q ~Uq ~�w  sq ~ 'D�Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_longst mount_longs:mxq ~9mq ~9lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9vsq ~ L�yT^uq ~ O   q ~ zt longsw  	�sq ~ 'N�s�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~3t nashua:nxq ~9~q ~9}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ L�A�uq ~ O   q ~3w  	 sq ~ '�\)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ L׺$�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�w'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_forakert mount_foraker:mxq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ L���uq ~ O   q ~ zt forakerw  sq ~ 'Oڒsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt south_gate_cat south_gate_ca:cxq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ LE�\�uq ~ O   q ~ Qq ~ �q ~
�t gatew  �sq ~ '�-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
appleton:nxq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ LFLG�uq ~ O   q ~�w  fsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fort_lauderdale_flt fort_lauderdale_fl:cxq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ L�8yvuq ~ O   q ~ Qq ~ �q ~ �t 
lauderdalew  �sq ~ '͊�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t north_little_rockt north_little_rock:nxq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ L���ruq ~ O   q ~Uq ~�q ~�w  sq ~ 'Y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~9�sq ~ L�$9ruq ~ O   q ~ Qq ~#q ~ �w   �sq ~ '~cBLsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_north_palisadet mount_north_palisade:mxq ~9�q ~9�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:sq ~ LH%�ouq ~ O   q ~ zq ~Ut palisadew  �sq ~ '�v�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~:
q ~:	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:sq ~ L����uq ~ O   q ~Nq ~q ~w  �sq ~ 'I�4�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t st_pault 	st_paul:nxq ~:q ~:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~: sq ~ L 6%�uq ~ O   q ~Nq ~
�w  �sq ~ '�~�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*Axq ~:'q ~:&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:-sq ~ LI�v*uq ~ O   q ~�w  	sq ~ '>�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~:4q ~:3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~::sq ~ LS�F$uq ~ O   q ~�q ~�q ~ �w  �sq ~ '_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~:Aq ~:@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:Gsq ~ L�W�uq ~ O   q ~ Qq ~ �q ~Ww  usq ~ '�-r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~_xq ~:Nq ~:Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:Tsq ~ L8�yuq ~ O   q ~ Qq ~ �q ~jw  �sq ~ '&`�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3�xq ~:[q ~:Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:asq ~ LS,��uq ~ O   q ~�q ~(�w   �sq ~ '��msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#0xq ~:hq ~:gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:nsq ~ Lz���uq ~ O   q ~�w  �sq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)�xq ~:uq ~:tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:{sq ~ L�~�uq ~ O   q ~ �q ~)�q ~ �w  �sq ~ '7>�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L�;�Euq ~ O   q ~ Qq ~1�w  	Isq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L`��uq ~ O   q ~�q ~uw  Usq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ LĴD�uq ~ O   q ~ Qq ~ �q ~�w  ~sq ~ '�~z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L���cuq ~ O   q ~ �q ~ �w  sq ~ '%W�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L�)�uq ~ O   q ~ gw  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!Ixq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L��guq ~ O   q ~ Qq ~ Rq ~ Sq ~fw  �sq ~ 'xe��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ Lp7Kuq ~ O   q ~�q ~�w  psq ~ '�
(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L���uq ~ O   q ~ Qq ~ �q ~ Rw  �sq ~ '4Y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L�eSuq ~ O   q ~�q ~5w   �sq ~ '�2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~:�q ~:�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:�sq ~ L!�|uq ~ O   q ~�q ~�w  sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~;q ~;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;
sq ~ L�Nuq ~ O   q ~�w  sq ~ 'f�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	wichita:nxq ~;q ~;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;sq ~ LO�Z�uq ~ O   q ~�w  �sq ~ 'w�Iq ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~;q ~;sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~;#sq ~ L 4dOuq ~ O   t passw  
<sq ~ 'q�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~2t minneapolis:nxq ~;+q ~;*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;3sq ~ LzbQ}uq ~ O   q ~2w  Hsq ~ '8���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt simi_valley_cat simi_valley_ca:cxq ~;:q ~;9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;Csq ~ L�{Ouq ~ O   t simiq ~q ~ �w  �sq ~ '=���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~,�t 
glendale:nxq ~;Kq ~;Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;Ssq ~ L�P�Buq ~ O   q ~,�w  �sq ~ '
��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~;Zq ~;Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;`sq ~ LӴ�*uq ~ O   q ~�q ~�w  �sq ~ '��Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~;gq ~;fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;msq ~ L��3>uq ~ O   q ~ Qq ~ �q ~2�w  sq ~ '��Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~;tq ~;ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;zsq ~ LKc�[uq ~ O   q ~�q ~�q ~Fw  sq ~ '�Osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L%���uq ~ O   q ~ Qq ~'�q ~ �w  	sq ~ '���bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L5{Duq ~ O   q ~ Qq ~ �q ~�w  sq ~ '  ��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~;�q ~w  	�sq ~ 'Uo�|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt rockford_ilt rockford_il:cxq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L�U�Duq ~ O   q ~ Qq ~ �q ~3sw  	Ksq ~ '#�6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
cranston:nxq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ Lfd�uq ~ O   q ~�w  �sq ~ '9{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L�_�fuq ~ O   q ~	�q ~�w  ssq ~ '��M�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L{�uq ~ O   q ~ Qq ~ Rq ~ Sq ~+Vw  lsq ~ 'E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ Lz���uq ~ O   q ~ Qq ~*q ~ �w  sq ~ '��#Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L���uq ~ O   q ~ �q ~ �q ~"w   {sq ~ 'WA��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~;�q ~;�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~;�sq ~ L+��uq ~ O   q ~Fq ~"w  sq ~ '�`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~<q ~< sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<sq ~ L���uq ~ O   q ~�q ~#w  sq ~ 'ĥS�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~<q ~<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<sq ~ ḶP�uq ~ O   q ~-�q ~#w  �sq ~ '{Le�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2xq ~<q ~<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<!sq ~ L
I��uq ~ O   q ~ Qq ~ �q ~ zq ~�w  Asq ~ '4,K[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~<(q ~<'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<.sq ~ L�Wҧuq ~ O   q ~Tq ~�w  jsq ~ '�C��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~<5q ~<4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<;sq ~ L�,�]uq ~ O   q ~Uq ~�q ~�q ~ �w   �sq ~ '�S�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~<Csq ~ L�ۂuq ~ O   t totalw  
&sq ~ 'bECsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~3t minnesota:sxq ~<Kq ~<Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<Ssq ~ L����uq ~ O   q ~ Qq ~ Rq ~ Sq ~3w  �sq ~ '�Jysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t 	bristol:nxq ~<Zq ~<Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<bsq ~ L���uq ~ O   q ~w  �sq ~ '�t�vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	skokie_ilt skokie_il:cxq ~<iq ~<hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<rsq ~ L�U6�uq ~ O   q ~"Nw  �sq ~ 'e��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6xq ~<yq ~<xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<sq ~ L�uq ~ O   q ~
/q ~#w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L��R�uq ~ O   q ~/q ~0w  csq ~ '���{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	toledo_oht toledo_oh:cxq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L��0�uq ~ O   t toledoq ~	�w  Psq ~ '�z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ LɛE�uq ~ O   q ~gq ~hw  �sq ~ 'ؤ�asq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	lorain_oht lorain_oh:cxq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L3�uq ~ O   q ~�q ~�w  Tsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L�y�uq ~ O   q ~ Qq ~ �q ~�q ~�w   �sq ~ '�R�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L,v��uq ~ O   q ~&�q ~�w  'sq ~ 'հ-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ Lg(Nuq ~ O   q ~�q ~w  �sq ~ 'p�*�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L�	Y�uq ~ O   q ~�q ~ �w  �sq ~ '��_sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0�xq ~<�q ~<�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~<�sq ~ L����uq ~ O   q ~ Qq ~ �q ~0�w  �sq ~ '�|a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt west_palm_beach_flt west_palm_beach_fl:cxq ~=q ~=sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=sq ~ L����uq ~ O   q ~ Qq ~ �q ~t palmq ~	bw  sq ~ '/�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt west_covina_cat west_covina_ca:cxq ~=q ~=sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=sq ~ L0�f}uq ~ O   q ~ Qq ~ �q ~t covinaw  �sq ~ '�n2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$oxq ~=$q ~=#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=*sq ~ Lc�
uq ~ O   q ~ �q ~$zw  	Vsq ~ '���xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t cincinnati:nxq ~=1q ~=0sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=9sq ~ L��uq ~ O   q ~�w   �sq ~ '�33�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;;xq ~=@q ~=?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=Fsq ~ LPAguq ~ O   q ~ Qq ~ �q ~;Fq ~w   �sq ~ '}X�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t livoniat 	livonia:nxq ~=Mq ~=Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=Vsq ~ L ͎uq ~ O   q ~=Ow  	�sq ~ '�4Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<jxq ~=]q ~=\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=csq ~ L+�uq ~ O   q ~"Nq ~Uw  	sq ~ 'I �q ~�sq ~ sq ~ sq ~ 
w   q ~Aq ~1vxq ~=iq ~=hsq ~ @q ~�sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~=mq ~�w   Fsq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~-�t pueblo:nxq ~=rq ~=qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=zsq ~ Lž�uq ~ O   q ~-�w  	sq ~ '<}�Osq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t chula_vistat chula_vista:nxq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L��t�uq ~ O   t chulat vistaw  sq ~ '�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt gainesville_flt gainesville_fl:cxq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L�A�Auq ~ O   t gainesvilleq ~�w  	psq ~ '�6q�q ~�sq ~ sq ~ sq ~ J   w   q ~5xq ~=�q ~=�sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~=�sq ~ L 5�?uq ~ O   q ~6w  	�sq ~ 'v��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L���uq ~ O   q ~ Rq ~ Sq ~�w  �sq ~ 'J �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ Lk�cUuq ~ O   q ~$�q ~	bq ~ �w  �sq ~ 'P��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	daly_cityt daly_city:nxq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L݇�uq ~ O   q ~�q ~ �w  	/sq ~ '��M2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L��W�uq ~ O   q ~ Rq ~ Sq ~w  sq ~ '��Nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<�xq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L����uq ~ O   q ~�w  Isq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#0xq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~=�sq ~ L�� �uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�i';sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~=�q ~=�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>sq ~ L\��uq ~ O   q ~)q ~Aw  �sq ~ 'D"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt middletown_njt middletown_nj:cxq ~>q ~>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>sq ~ LA��uq ~ O   t 
middletownq ~(�w  sq ~ 'ޠ�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~>q ~>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>#sq ~ L��c�uq ~ O   q ~ Qq ~ �q ~Uq ~�w  �sq ~ 'B��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_wrangellt mount_wrangell:mxq ~>*q ~>)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>3sq ~ LDJuq ~ O   q ~ zt wrangellw  �sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt cheektowaga_nyt cheektowaga_ny:cxq ~>;q ~>:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>Dsq ~ L~*+fuq ~ O   q ~*q ~�w  �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~gt idaho:nxq ~>Kq ~>Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>Ssq ~ L��kuq ~ O   q ~gw  \sq ~ '*��Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Yxq ~>Zq ~>Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>`sq ~ L*�_uq ~ O   q ~ Qq ~ �q ~ fw  }sq ~ '/y[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~>gq ~>fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>msq ~ L*�uq ~ O   q ~1q ~�w  �sq ~ 'N|�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~>usq ~ LN{��uq ~ O   t whitneyw  
*sq ~ '�Ղ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~>}q ~>|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~�xq ~>�sq ~ L 3�uq ~ O   t doq ~ w   !sq ~ '-�'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
buffalo_nyt buffalo_ny:cxq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>�sq ~ L�Uuq ~ O   q ~ Qq ~ �q ~�w   �sq ~ '�z[#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t allegheny_rivert allegheny_river:rxq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>�sq ~ L��GAuq ~ O   t 	alleghenyq ~ �w  �sq ~ '�<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0xq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>�sq ~ L��.uq ~ O   q ~ q ~;w  �sq ~ '<\�q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~>�q ~>�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~>�sq ~ Lī��uq ~ O   t passesw  	�sq ~ ' 6�$sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~>�sq ~ L 6M�uq ~ O   q ~*w   sq ~ 'Ċ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>�sq ~ Ljh�luq ~ O   q ~�q ~�w  �sq ~ '	�,Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t ogden:nxq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>�sq ~ LL�suq ~ O   q ~�w  {sq ~ '9{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>�sq ~ L?7�!uq ~ O   q ~�q ~Tw  osq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~>�q ~>�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~? sq ~ LO��uq ~ O   q ~�q ~�q ~ w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~?q ~?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?sq ~ L1?�uq ~ O   q ~ �w  1sq ~ '�2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~?q ~?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?sq ~ L_�duq ~ O   q ~�w  $sq ~ 'Y\�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7�xq ~?!q ~? sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?'sq ~ L!H&1uq ~ O   q ~7�q ~5w  3sq ~ '��\nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~?.q ~?-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?4sq ~ Lz-�uq ~ O   q ~ Qq ~ �q ~.�w  
sq ~ 'z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~?;q ~?:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?Asq ~ L�$��uq ~ O   q ~�q ~�q ~�w  vsq ~ '��<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~?Hq ~?Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?Nsq ~ L�E�(uq ~ O   q ~ Qq ~�w  �sq ~ '�oZq ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~?Tq ~?Ssq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~?Xsq ~ L �uq ~ O   t forw  	�sq ~ '�(Ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt chattanooga_tnt chattanooga_tn:cxq ~?`q ~?_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?isq ~ L'uq ~ O   q ~ Qq ~ �q ~8�w  �sq ~ '���lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'Pxq ~?pq ~?osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?vsq ~ L)Ac�uq ~ O   q ~'[w  0sq ~ 'F=zOsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.Lxq ~?}q ~?|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L�۫Fuq ~ O   q ~.Wq ~�q ~�w  �sq ~ 'gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L�W{uq ~ O   q ~"q ~ �w  �sq ~ '�Z�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L>6��uq ~ O   q ~q ~ �q ~w  sq ~ '�v�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~jt 	chicago:nxq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L,w�uq ~ O   q ~jw  3sq ~ '`�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	kendall:nxq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L��COuq ~ O   q ~�w  �sq ~ '�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt waukegan_ilt waukegan_il:cxq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L1�۴uq ~ O   t waukeganq ~5w  sq ~ '玘Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t irvingt irving:nxq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L����uq ~ O   q ~?�w  'sq ~ '	��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ L�U,�uq ~ O   q ~Uq ~�t scw  �sq ~ '��y+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~?�sq ~ LJ�8uq ~ O   q ~!�q ~ gw  Nsq ~ '`
�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~)?t 	dubuque:nxq ~?�q ~?�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@sq ~ Lw2�uq ~ O   q ~)?w  �sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3xq ~@q ~@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@sq ~ L��uq ~ O   q ~~w  �sq ~ '�P��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t huntington_beacht huntington_beach:nxq ~@q ~@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@#sq ~ Lc��?uq ~ O   q ~�q ~	bw  �sq ~ '�;L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt parma_oht 
parma_oh:cxq ~@*q ~@)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@3sq ~ LX3uq ~ O   q ~�w  :sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~@:q ~@9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@@sq ~ L�^iuq ~ O   q ~ Qq ~ �q ~'w  �sq ~ '2"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Kxq ~@Gq ~@Fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@Msq ~ L̈��uq ~ O   q ~ Qq ~ �q ~Vw  dsq ~ '�D��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~-Yt woodbridge:nxq ~@Tq ~@Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@\sq ~ L:��uq ~ O   q ~-Yw  �sq ~ 'a6_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~@cq ~@bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@isq ~ LѦ��uq ~ O   q ~ Qq ~ �q ~+�w  �sq ~ 'J��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
/t 
lakewood:nxq ~@pq ~@osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@xsq ~ L����uq ~ O   q ~
/w  .sq ~ '�k �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
west_allist west_allis:nxq ~@q ~@~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ LF:�uq ~ O   q ~q ~ww  �sq ~ '�B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~@�sq ~ L��[uq ~ O   t whichw   sq ~ 'M���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,�xq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ Ln`�uq ~ O   q ~ Qq ~ �q ~(�w   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ L���uq ~ O   q ~�w  Tsq ~ '4��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~@�sq ~ L4<Wuq ~ O   q ~ zw  
)sq ~ '�[=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ L�n��uq ~ O   q ~�q ~	�w  �sq ~ 'ZS߲sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt largo_flt 
largo_fl:cxq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ L�0Juq ~ O   t largoq ~"w  Asq ~ '��V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ LU���uq ~ O   q ~w  �sq ~ '�i sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.Lxq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~@�sq ~ LsOuq ~ O   q ~.Ww  �sq ~ 'Sz�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt green_bay_wit green_bay_wi:cxq ~@�q ~@�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A sq ~ L
��uq ~ O   q ~q ~#q ~xw  �sq ~ 'x��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Aq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Asq ~ L��uq ~ O   q ~'w  �sq ~ 'w�isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~Aq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~Asq ~ L  uq ~ O   q ~ Sw   >sq ~ 'wK-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
anaheim_cat anaheim_ca:cxq ~A!q ~A sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A*sq ~ Lر�Yuq ~ O   q ~ Qq ~ �t anaheimw  	9sq ~ '�G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~A2q ~A1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A8sq ~ Lw$Тuq ~ O   q ~&q ~Tw  sq ~ 'x��>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt metairie_lat metairie_la:cxq ~A?q ~A>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~AHsq ~ L�hp.uq ~ O   q ~ Qq ~ �t metairiew  isq ~ '�dRsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~APq ~AOsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~AVsq ~ L�fnxuq ~ O   q ~�q ~"w  Dsq ~ '�S��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5cxq ~A]q ~A\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Acsq ~ LY�r|uq ~ O   q ~ Qq ~�w  �sq ~ 'd���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~Ajq ~Aisq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Apsq ~ L��
�uq ~ O   q ~ Qq ~ �q ~$�q ~	bw  'sq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Awq ~Avsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A}sq ~ L��yuq ~ O   q ~�q ~ �q ~ �w   �sq ~ '�.��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ut euclid:nxq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L���2uq ~ O   q ~Uw  isq ~ '�Wusq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t dayton:nxq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L�4Huuq ~ O   q ~�w  	sq ~ '� G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L2�R(uq ~ O   q ~w  wsq ~ '_��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	camden_njt camden_nj:cxq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L�y�uq ~ O   q ~#w   �sq ~ '!�&�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
jackson_mst jackson_ms:cxq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L����uq ~ O   q ~Ut msw  �sq ~ '��asq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt pasadena_cat pasadena_ca:cxq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ LG�J�uq ~ O   q ~w  �sq ~ 'ТY�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\xq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L�OUuq ~ O   q ~�q ~4q ~ Rw  �sq ~ '
�)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~t hawaii:sxq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~A�sq ~ L0S��uq ~ O   q ~q ~ Rw  �sq ~ '�&��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>�xq ~A�q ~A�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Bsq ~ L�E�Zuq ~ O   q ~�q ~�w  	(sq ~ '`j.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
high_pointt high_point:nxq ~B	q ~Bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Bsq ~ LI0uq ~ O   q ~�q ~�w  sq ~ '6�`�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)4xq ~Bq ~Bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Bsq ~ Lo@�Suq ~ O   q ~)?q ~�w  �sq ~ ' *!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*oxq ~B&q ~B%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B,sq ~ L����uq ~ O   q ~*zw  	sq ~ '��z�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~B4sq ~ L��luq ~ O   t 	guadalupew  
sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~B<q ~B;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~BBsq ~ L�*�Tuq ~ O   q ~�q ~�w  sq ~ '�j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~BIq ~BHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~BOsq ~ L���uq ~ O   q ~�q ~ �w  =sq ~ '���Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~BVq ~BUsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B\sq ~ L�&(�uq ~ O   q ~�q ~�q ~ gw  vsq ~ '���Gq ~�sq ~ sq ~ sq ~ J   w   q ~Mq ~"exq ~Bbq ~Basq ~ @q ~�sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~Bfsq ~ L��3uq ~ O   q ~?w  
\sq ~ '��_sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	racine_wit racine_wi:cxq ~Bmq ~Blsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Bvsq ~ L���uq ~ O   q ~�w  ssq ~ '|W��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~B}q ~B|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ LjU�/uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w   �sq ~ 'X@?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'?xq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ L8�0�uq ~ O   q ~'Jw  �sq ~ 'J�7Asq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~t north_dakota:sxq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ L�a�uq ~ O   q ~ Rq ~ Sq ~Uq ~
�w  	�sq ~ '��ژsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~	!xq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~B�sq ~ L��7,uq ~ O   q ~5�w   Isq ~ 'Ǟ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt colorado_springs_cot colorado_springs_co:cxq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ Ly�B�uq ~ O   q ~ Qq ~ �q ~#t springsw   �sq ~ '�y�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt tempe_azt 
tempe_az:cxq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ L˴�(uq ~ O   t tempeq ~pw  �sq ~ '�(��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ L0��quq ~ O   q ~�w  	�sq ~ '�K��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~mxq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ L��\�uq ~ O   q ~�t arizonaw  7sq ~ '$UXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t indianapolist indianapolis:nxq ~B�q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~B�sq ~ L"E�uq ~ O   q ~B�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Txq ~C q ~B�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Csq ~ LF�uq ~ O   q ~ q ~=q ~ �w  �sq ~ '�&�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt chula_vista_cat chula_vista_ca:cxq ~Cq ~Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Csq ~ L�~0�uq ~ O   q ~=�q ~=�q ~ �w  �sq ~ '˸��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~Cq ~Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C#sq ~ L�葉uq ~ O   q ~ Qq ~8�q ~ �w  	sq ~ '�Q�Osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~C*q ~C)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C0sq ~ L 9uq ~ O   q ~hq ~ Sq ~�w  'sq ~ 'q�j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
fort_wortht fort_worth:nxq ~C7q ~C6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C@sq ~ L��uq ~ O   q ~ �t worthw  �sq ~ '4��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~CHq ~CGsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~CNsq ~ Lf9z�uq ~ O   q ~�q ~�w  �sq ~ '$,�Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~04xq ~CUq ~CTsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C[sq ~ L�
�uq ~ O   q ~0?q ~Uw  �sq ~ '?�3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~Cbq ~Casq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Chsq ~ LQ�k�uq ~ O   q ~fw   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Coq ~Cnsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Cusq ~ Ll��/uq ~ O   q ~�q ~=w  �sq ~ 'X�'$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~C|q ~C{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ L[7�uq ~ O   q ~ q ~	bq ~=w   �sq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%�xq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ LK��Nuq ~ O   q ~ Qq ~ �q ~%5w  sq ~ '�O�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~!�t 	saginaw:nxq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ Lnϋ�uq ~ O   q ~!�w  sq ~ '��Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'xq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ LK���uq ~ O   q ~'q ~Uq ~�w  )sq ~ '�ƫsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ L� ��uq ~ O   q ~ Qq ~ �q ~�q ~�w  nsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8-xq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ L�}5�uq ~ O   q ~ Qq ~ �q ~�q ~�w  Dsq ~ 'ס,�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~wt schenectady:nxq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ L���uq ~ O   q ~ww  �sq ~ '9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t mesa:nxq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ L 3$uq ~ O   q ~�w  �sq ~ '"/�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t scotts_valleyt scotts_valley:nxq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~C�sq ~ LA��Kuq ~ O   q ~nq ~w  �sq ~ '��Q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~C�q ~C�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D sq ~ Lz���uq ~ O   q ~�w  �sq ~ '�W�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	duluth_mnt duluth_mn:cxq ~Dq ~Dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Dsq ~ L�H:uq ~ O   q ~�w  �sq ~ '
���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Dq ~Dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Dsq ~ L[���uq ~ O   q ~�w   �sq ~ '۫��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~D$q ~D#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D*sq ~ L)Bӵuq ~ O   q ~�w  �sq ~ '� 48sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t pennsylvania:nxq ~D1q ~D0sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D9sq ~ L2�R(uq ~ O   q ~w  �sq ~ ',8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~D@q ~D?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~DFsq ~ Lڄ�uq ~ O   q ~#w  ?sq ~ '��5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%Qxq ~DMq ~DLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~DSsq ~ L�Ŗquq ~ O   q ~ Qq ~ �q ~%\w  ksq ~ 'V��fq ~�sq ~ sq ~ sq ~ J   w   q ~�q ~�xq ~DYq ~DXsq ~ @q ~�sq ~ Go��    sq ~ sq ~ J   w   q ~q ~xq ~D]q ~&�w  
>sq ~ '��DGsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_uncompahgret mount_uncompahgre:mxq ~Dbq ~Dasq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Dksq ~ Lp.�uq ~ O   q ~ zt uncompahgrew  sq ~ '��(q ~�sq ~ sq ~ sq ~ J   w   q ~	!xq ~Drq ~Dqsq ~ @q ~�sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~Dvsq ~ L 3�uq ~ O   q ~3w  	�sq ~ 'E6��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t colorado_springst colorado_springs:nxq ~D}q ~D|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L���uq ~ O   q ~#q ~B�w  usq ~ '�U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!exq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L����uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�:68sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~2�t levittown:nxq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L����uq ~ O   q ~2�w  Gsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0�xq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L�N�Huq ~ O   q ~0�w  sq ~ 'p���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L��1uq ~ O   q ~fq ~ gw  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Hxq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ Lx�Fuq ~ O   q ~ Qq ~ �q ~Sw  �sq ~ 'Z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt thousand_oaks_cat thousand_oaks_ca:cxq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L���uq ~ O   q ~ Qq ~ �t thousandt oaksw  $sq ~ '�eP^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ L"V�uq ~ O   q ~ �q ~		w  �sq ~ 'c��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!exq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~D�sq ~ LS���uq ~ O   q ~�q ~w  6sq ~ '��[xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~	�t 
columbus:nxq ~D�q ~D�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Esq ~ L��7�uq ~ O   q ~	�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_kit_carsont mount_kit_carson:mxq ~Eq ~E
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Esq ~ L�ćuq ~ O   q ~ zt kitq ~*w  �sq ~ '��q ~�sq ~ sq ~ sq ~ J   w   q ~xq ~Eq ~Esq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~Esq ~ Ld�wuq ~ O   t populationsw  	�sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t mcallent 	mcallen:nxq ~E'q ~E&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E0sq ~ L4��ruq ~ O   q ~E)w   �sq ~ 'Q�l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~E7q ~E6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E=sq ~ L��uq ~ O   q ~ Qq ~ �q ~3q ~'�w  /sq ~ ' 4pq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~EEsq ~ L 3�1uq ~ O   t nextw  	�sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_crestone_needlet mount_crestone_needle:mxq ~EMq ~ELsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~EVsq ~ LM�4wuq ~ O   q ~ zt crestonet needlew  �sq ~ '�,�@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~~xq ~E_q ~E^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Eesq ~ L�#xuq ~ O   q ~�q ~�w  �sq ~ '�
�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bnxq ~Elq ~Eksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ersq ~ L�Fg�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '6���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~:xq ~Eyq ~Exsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Esq ~ LȇH%uq ~ O   t riversw   Vsq ~ '�Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t tahoet tahoe:lxq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L���uq ~ O   q ~q ~E�w  	
sq ~ 'ʃP sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L�gˏuq ~ O   q ~Uq ~ �w   zsq ~ '{g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ �^��tt <<e,t>,<<e,i>,i>>q ~ �sq ~ �H���t 	<<e,i>,i>q ~Jq ~t sumt sum:<<e,t>,<<e,i>,i>>xq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~E�sq ~ L�ۂuq ~ O   q ~<Fw   /sq ~ '�zxgsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L�s��uq ~ O   q ~Nq ~ �w  �sq ~ 'O��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L?-��uq ~ O   q ~�q ~�q ~ �w  �sq ~ 'Y���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@�xq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L��uq ~ O   q ~q ~#q ~*w  �sq ~ '"��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L�{��uq ~ O   q ~ Qq ~ �q ~+�w  �sq ~ '��Ԙsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	vermont:nxq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~E�sq ~ L�yIuq ~ O   q ~�w   �sq ~ '�?Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~E�q ~E�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Fsq ~ L�z`�uq ~ O   q ~B�q ~B�w  �sq ~ ' 0�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~Fq ~Fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~Fsq ~ L 0R/uq ~ O   q ~`q ~*�w   6sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~Fq ~Fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Fsq ~ L�z!uq ~ O   q ~w  	�sq ~ '�e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt pittsburgh_pat pittsburgh_pa:cxq ~F"q ~F!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F+sq ~ L�gj�uq ~ O   t 
pittsburghw  	ysq ~ '{-M�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~{xq ~F3q ~F2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F9sq ~ Lj�,uq ~ O   q ~ Qq ~ �q ~�w  Csq ~ '�ޑ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~F@q ~F?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~FFsq ~ L��uq ~ O   q ~Uq ~ �q ~�w  	Bsq ~ '-��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5�xq ~FMq ~FLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~FSsq ~ L���uq ~ O   q ~Iw  �sq ~ 'U!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#yxq ~FZq ~FYsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F`sq ~ L�&uq ~ O   q ~�q ~#�w  �sq ~ 't�(Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~1Ct winston-salem:nxq ~Fgq ~Ffsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Fosq ~ L�uq ~ O   q ~1Cw   sq ~ '#<߮sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Fvq ~Fusq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F|sq ~ L�3O�uq ~ O   q ~q ~ �w  �sq ~ 'EX�zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ LE=g�uq ~ O   q ~ Qq ~ �q ~Uq ~ �w  +sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ L���uq ~ O   q ~ Qq ~ �q ~�w  4sq ~ 'i�Euq ~=sq ~ sq ~ sq ~ 
w   q ~Hxq ~F�q ~F�sq ~ @q ~Lsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~F�q ~Qw   'sq ~ 'PLsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ LDp�uq ~ O   q ~ Qq ~ �q ~gq ~hw  nsq ~ '�ӏ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~?�xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ L�s�uq ~ O   q ~?�q ~Uw  9sq ~ '�oRsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ LaF��uq ~ O   q ~ Rq ~ Sq ~"w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ L؛��uq ~ O   q ~q ~Uw  sq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ L6�uq ~ O   q ~ Qq ~ �q ~Nq ~�w  �sq ~ '��dCsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ L}2'buq ~ O   q ~ Qq ~ Rq ~ Sq ~Wq ~ Sq ~Xw  �sq ~ '�{%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~F�q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~F�sq ~ L�~��uq ~ O   q ~�q ~ Rw  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_belfordt mount_belford:mxq ~G q ~F�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G	sq ~ L��g�uq ~ O   q ~ zt belfordw  fsq ~ '���[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	lowell_mat lowell_ma:cxq ~Gq ~Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Gsq ~ LGv�uq ~ O   t lowellq ~�w  sq ~ '0�90sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt mesquite_txt mesquite_tx:cxq ~G"q ~G!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G+sq ~ L�n��uq ~ O   t mesquiteq ~ �w  �sq ~ 'Տ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Dxq ~G3q ~G2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G9sq ~ L���ruq ~ O   q ~ Qq ~ �q ~�w  sq ~ 'XF��q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~G?q ~G>sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~GCsq ~ L�7auq ~ O   q ~�w  
sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~GJq ~GIsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~GPsq ~ L�nӫuq ~ O   q ~
Yq ~"w  �sq ~ 'l~^�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A@xq ~GWq ~GVsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G]sq ~ L�/��uq ~ O   q ~AKw  	isq ~ 'n�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~Gdq ~Gcsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Gjsq ~ L�t�uq ~ O   q ~,q ~ �w  sq ~ 's�D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Gqq ~Gpsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Gwsq ~ L���uq ~ O   q ~�q ~"w  `sq ~ '�f��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t north_platte_rivert north_platte_river:rxq ~G~q ~G}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L��>*uq ~ O   q ~ Qq ~Uq ~5w  �sq ~ '��}asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<�xq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L�+�uq ~ O   q ~<�q ~�w  �sq ~ '�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~?�t 
waukegan:nxq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L"��muq ~ O   q ~?�w  �sq ~ '3|�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L�jO�uq ~ O   q ~ Qq ~ �q ~Fw  �sq ~ 'g"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L���5uq ~ O   q ~+q ~�q ~�w   �sq ~ '9#��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'0t 	ontario:nxq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L�=Juq ~ O   q ~'0w  wsq ~ '�-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=�xq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L˚�Xuq ~ O   q ~=�q ~"w  Qsq ~ '<F��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt huntington_wvt huntington_wv:cxq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L]uq ~ O   q ~�q ~�w  �sq ~ '%Z	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~G�sq ~ L	��Vuq ~ O   q ~ Rq ~ Sq ~�q ~Fw  �sq ~ '?Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(#xq ~G�q ~G�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Hsq ~ L�|5quq ~ O   q ~(.w  sq ~ 'o�S�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~7�t warren:nxq ~H
q ~H	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Hsq ~ LН$�uq ~ O   q ~7�w  Tsq ~ 'B���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t santa_barbarat santa_barbara:nxq ~Hq ~Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H"sq ~ L��<tuq ~ O   q ~ q ~5w  �sq ~ '��� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'rxq ~H)q ~H(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H/sq ~ Lh-uq ~ O   q ~ Qq ~ �q ~'}w  sq ~ 'ٙ}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~H6q ~H5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H<sq ~ L����uq ~ O   q ~)q ~)q ~w  sq ~ 'I7Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;�xq ~HCq ~HBsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~HIsq ~ L�Q�uq ~ O   q ~3sw  Lsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~HPq ~HOsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~HVsq ~ L�L�uq ~ O   q ~�q ~ �w  �sq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~H]q ~H\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Hcsq ~ L-�
uq ~ O   q ~ >w  �sq ~ ' 6�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Hksq ~ L 6M�uq ~ O   q ~Tw  	�sq ~ '1�{q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Hssq ~ L1_<uq ~ O   t milesw  	�sq ~ '�?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~H{q ~Hzsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L�V�uq ~ O   q ~ �q ~ �w  asq ~ 'H<�usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L���7uq ~ O   q ~�q ~"w  osq ~ '�4��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~0?t 
evanston:nxq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L	�9�uq ~ O   q ~0?w  sq ~ '�l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L g�Wuq ~ O   q ~ �q ~Nw  �sq ~ '- 8[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0xq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L��Ruq ~ O   q ~;q ~~w  	dsq ~ 'ȗ
Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t cicero:nxq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L����uq ~ O   q ~w  =sq ~ '�&sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!uxq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L:�{uq ~ O   q ~ �q ~!�w  �sq ~ '
TR�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~wt lawton:nxq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L��$�uq ~ O   q ~ww  sq ~ '? ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/4xq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ Lʸ�>uq ~ O   q ~
�q ~�w  �sq ~ 'wg��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~H�q ~H�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~H�sq ~ L��uq ~ O   q ~q ~q ~ �w  �sq ~ '�h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Iq ~Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I	sq ~ L4x>uq ~ O   q ~�q ~Uq ~�w  �sq ~ 'Er[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	topeka_kst topeka_ks:cxq ~Iq ~Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Isq ~ L��uq ~ O   q ~1�q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~I q ~Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I&sq ~ L�,e�uq ~ O   q ~�w  �sq ~ '.��0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~I-q ~I,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I3sq ~ L��uq ~ O   q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~I:q ~I9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I@sq ~ La��uq ~ O   q ~ Qq ~ �q ~�w  	�sq ~ '=�a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0Uxq ~IGq ~IFsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~IMsq ~ L{A�iuq ~ O   q ~ Qq ~ �q ~�q ~�w  �sq ~ '<h��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt charleston_sct charleston_sc:cxq ~ITq ~ISsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I]sq ~ L]�uq ~ O   q ~�w  �sq ~ 'd1Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~Idq ~Icsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ijsq ~ LíQ�uq ~ O   q ~Dq ~w  Ysq ~ '�A�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
pontiac_mit pontiac_mi:cxq ~Iqq ~Ipsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Izsq ~ L$�Ruq ~ O   t pontiacq ~Tw  �sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t san_leandrot san_leandro:nxq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ L:�{uq ~ O   q ~ �q ~!�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt springfield_mat springfield_ma:cxq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ L��Iuq ~ O   q ~Fq ~�w  9sq ~ 'm6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t townt town:<lo,t>xq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~I�sq ~ L��_uq ~ O   t townsw   7sq ~ '�-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ LO>�uq ~ O   q ~ Rq ~ Sq ~�q ~�w  �sq ~ '?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ L����uq ~ O   q ~ Qq ~ �q ~Uw  sq ~ '>ޕ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t lynchburg:nxq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ L#�uq ~ O   q ~�w  !sq ~ ' �~;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt savannah_gat savannah_ga:cxq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ L���uq ~ O   t savannahq ~+w   �sq ~ '7�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~St 	wyoming:sxq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~I�sq ~ L��uq ~ O   q ~Sq ~ Rw  Gsq ~ 'zO	>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"�xq ~I�q ~I�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ L��i`uq ~ O   q ~ Qq ~ �q ~
/w  -sq ~ '�	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9�xq ~J	q ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ L�ψuq ~ O   q ~ �q ~9�q ~�w  	�sq ~ 'S4�Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Jq ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jsq ~ LўfYuq ~ O   q ~�q ~�w  sq ~ '��q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~J#q ~J"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J)sq ~ L�}Suq ~ O   q ~q ~=q ~"w  �sq ~ '�Z�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~><xq ~J0q ~J/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J6sq ~ L5�C#uq ~ O   q ~*w  �sq ~ '| �{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8^xq ~J=q ~J<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~JCsq ~ L /��uq ~ O   q ~8iq ~/Lw   �sq ~ '�=:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~}xq ~JJq ~JIsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~JPsq ~ L�DWIuq ~ O   q ~�q ~�q ~uw  �sq ~ '�b8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~"t clearwater:nxq ~JWq ~JVsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J_sq ~ L՛�(uq ~ O   q ~"w  �sq ~ '[��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(xq ~Jfq ~Jesq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Jlsq ~ L�δuq ~ O   q ~3q ~	bq ~"w  sq ~ '  ��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Jtsq ~ L  iuq ~ O   t itw  
3sq ~ '2){�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt independence_mot independence_mo:cxq ~J|q ~J{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L,���uq ~ O   q ~ Qq ~ �q ~gw  �sq ~ 'Aj �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A"xq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L�Т�uq ~ O   q ~A-q ~"w  �sq ~ '6�H�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t dakota_rivert dakota_river:rxq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L�d*]uq ~ O   q ~ Qq ~
�w  [sq ~ '&\��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~-�t oxnard:nxq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L�8l�uq ~ O   q ~-�w   sq ~ 'w=��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Axq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ LsVĶuq ~ O   q ~ Qq ~ �q ~Lw  	sq ~ 'H�b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L f�fuq ~ O   q ~ Qq ~�w  ^sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L]o�	uq ~ O   q ~�q ~!q ~"�w  sq ~ '4���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0xq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L���uq ~ O   q ~ Qq ~ �q ~;w  *sq ~ 'Mb�Asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6�xq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L���uq ~ O   q ~6�w  �sq ~ '(?��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*Pxq ~J�q ~J�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~J�sq ~ L���muq ~ O   q ~ Qq ~ �q ~*[q ~*\w  �sq ~ '��m{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Kq ~Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ksq ~ L2�{�uq ~ O   q ~q ~q ~ �q ~�w  sq ~ 'Y5�\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*Pxq ~Kq ~Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ksq ~ L���Guq ~ O   q ~*[q ~*\q ~Tw   �sq ~ '�cn�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~K q ~Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K&sq ~ Lp��uq ~ O   q ~3q ~'�q ~ w  sq ~ '��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t 
abingdon:nxq ~K-q ~K,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K5sq ~ LU���uq ~ O   q ~w  sq ~ '�)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~K<q ~K;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~KBsq ~ L���uq ~ O   q ~ Qq ~�q ~ �w   sq ~ '�"4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~KIq ~KHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~KOsq ~ L>i�uq ~ O   q ~ �q ~�w  �sq ~ '���"q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~KUq ~KTsq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~KYsq ~ L���uq ~ O   q ~ Rw  
Usq ~ '�J��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~K`q ~K_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Kfsq ~ LQ��uq ~ O   q ~�q ~ w  �sq ~ 'F_��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt glendale_cat glendale_ca:cxq ~Kmq ~Klsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Kvsq ~ L�P�Buq ~ O   q ~,�w  �sq ~ '}�UUsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~K}q ~K|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L��/�uq ~ O   q ~-�q ~"w  7sq ~ 'v�1�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t iowa:sxq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L 1j�uq ~ O   q ~�w   �sq ~ '�/>�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Xt tampa:nxq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L�e�uq ~ O   q ~Xw  �sq ~ 'e�-"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,�xq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L\uq ~ O   q ~,�q ~B�w  �sq ~ '8���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"sxq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L\S��uq ~ O   q ~�q ~#w  fsq ~ '"�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L�
�uq ~ O   q ~Fq ~5w  Wsq ~ 'e�$;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L����uq ~ O   q ~. q ~w  sq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L�cuq ~ O   q ~�q ~w  msq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(xq ~K�q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~K�sq ~ L�zHxuq ~ O   q ~ Qq ~ �q ~3w   lsq ~ '�\�pq ~�sq ~ sq ~ sq ~ J   w   q ~5xq ~K�q ~K�sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~K�sq ~ Lm\4�uq ~ O   q ~�w  
/sq ~ '�Ϥsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%�xq ~L q ~K�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Lsq ~ L�~Z�uq ~ O   q ~q ~w  sq ~ '��$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ht gary:nxq ~Lq ~Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Lsq ~ L 0L�uq ~ O   q ~hw  	�sq ~ '��L=sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~Lq ~Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L"sq ~ Lm��(uq ~ O   q ~ Qq ~ �q ~�w   �sq ~ '�8qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=�xq ~L)q ~L(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L/sq ~ L���uq ~ O   q ~ Qq ~ �q ~=�w  �sq ~ 'ǂ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$oxq ~L6q ~L5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L<sq ~ L�+�uq ~ O   q ~ �q ~$zq ~ �w  Wsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~LCq ~LBsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~LIsq ~ L�.?�uq ~ O   q ~%w  sq ~ '�A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"�xq ~LPq ~LOsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~LVsq ~ L5�7uq ~ O   q ~"�q ~ �w  	>sq ~ 'W��"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~L]q ~L\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Lcsq ~ L+���uq ~ O   q ~ Qq ~ �q ~�q ~Ew  �sq ~ 'y���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
$xq ~Ljq ~Lisq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Lpsq ~ L��i`uq ~ O   q ~ Qq ~ �q ~
/w  -sq ~ 'P�=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5xq ~Lwq ~Lvsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L}sq ~ L�b�buq ~ O   q ~ Qq ~
�q ~5w  �sq ~ 'i���q ~sq ~ sq ~ sq ~ 
w   q ~Hxq ~L�q ~L�sq ~ @q ~sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~L�q ~!w   ;sq ~ '<AL�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L��
uq ~ O   q ~�q ~!w  �sq ~ ')���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t arvada:nxq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L��Wuq ~ O   q ~�w  sq ~ 'ΰ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~2�t pawtucket:nxq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L�١|uq ~ O   q ~2�w  sq ~ '��hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t san_juan_rivert san_juan_river:rxq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L�uq ~ O   q ~ �t juanq ~ �w  �sq ~ 'Z�A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ LN0$�uq ~ O   q ~�w  �sq ~ 'c��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt philadelphia_pat philadelphia_pa:cxq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L,��5uq ~ O   q ~�q ~w  Msq ~ 'f`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_whitet mount_white:mxq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L�uq ~ O   q ~ zq ~Nw  sq ~ '�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt indianapolis_int indianapolis_in:cxq ~L�q ~L�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~L�sq ~ L"E�uq ~ O   q ~B�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Mq ~Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Msq ~ L� �?uq ~ O   q ~�q ~ �w  \sq ~ '0���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~Mq ~Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Msq ~ L���<uq ~ O   q ~�q ~�w   ssq ~ '	R�Isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7yxq ~Mq ~Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M%sq ~ L�ՕWuq ~ O   q ~ Qq ~ �q ~7�w  Fsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t el_montet 
el_monte:nxq ~M,q ~M+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M5sq ~ L5��uq ~ O   q ~ �q ~`w  �sq ~ '.B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
kenosha_wit kenosha_wi:cxq ~M<q ~M;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~MEsq ~ L�R�uq ~ O   t kenoshaq ~*w  �sq ~ '~���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t washita_rivert washita_river:rxq ~MMq ~MLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~MVsq ~ LCG_&uq ~ O   q ~ Qt washitaw  �sq ~ 'J��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt reno_nvt 	reno_nv:cxq ~M^q ~M]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Mgsq ~ L���uq ~ O   q ~�q ~�w  .sq ~ '獯�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~*zt irvine:nxq ~Mnq ~Mmsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Mvsq ~ L����uq ~ O   q ~*zw  |sq ~ 'e�0*sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)�xq ~M}q ~M|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ LH��uq ~ O   q ~ Qq ~ �q ~ �q ~)�w  �sq ~ 'm�K{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ Lё�0uq ~ O   q ~�q ~Tw  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ L��w�uq ~ O   q ~ Qq ~ �q ~I�w  0sq ~ '�V��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ L��luq ~ O   q ~�w  Dsq ~ '��θsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t utah:nxq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ L 6�Duq ~ O   q ~w  �sq ~ '�@2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Mxq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ L���Luq ~ O   q ~Xq ~"w  �sq ~ '��nQq ~=sq ~ sq ~ sq ~ 
w   q ~Hq ~Hxq ~M�q ~M�sq ~ @q ~Lsq ~ Go��    sq ~ sq ~ J   w   q ~q ~xq ~M�q ~Qw   4sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~?axq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~M�sq ~ L�X��uq ~ O   q ~8�w  Bsq ~ 'ZLi�q ~�sq ~ sq ~ sq ~ J   w   q ~;xq ~M�q ~M�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~M�sq ~ L���uq ~ O   q ~ Rw  
$sq ~ '�a��q ~�sq ~ sq ~ sq ~ J   w   q ~Hxq ~M�q ~M�sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~M�q ~+$w  	�sq ~ 'zn�q ~�sq ~ sq ~ sq ~ J   w   q ~Exq ~M�q ~M�sq ~ @q ~�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~M�sq ~ Luq ~ O   t greatestw  	�sq ~ '�a=sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~M�q ~M�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Nsq ~ L���uq ~ O   q ~ Qq ~ �q ~L�w  Xsq ~ '�"Dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Nq ~Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Nsq ~ L� }�uq ~ O   q ~�q ~ Rw  hsq ~ 'Ͽ�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t youngstown:nxq ~Nq ~Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N!sq ~ L����uq ~ O   q ~�w  +sq ~ '3b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3xq ~N(q ~N'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N.sq ~ L���uq ~ O   q ~ Qq ~ �q ~~w  �sq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~G�xq ~N5q ~N4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N;sq ~ L�?�Xuq ~ O   q ~�q ~q ~ w  �sq ~ '��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t washington:nxq ~NBq ~NAsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~NJsq ~ L�,e�uq ~ O   q ~�w  �sq ~ 'C?Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0�xq ~NQq ~NPsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~NWsq ~ L�R�uq ~ O   q ~ Rq ~ Sq ~ w  	�sq ~ 'C�L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~N^q ~N]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ndsq ~ L�J��uq ~ O   q ~w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~pt charlotte:nxq ~Nkq ~Njsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Nssq ~ L]�4*uq ~ O   q ~pw  -sq ~ 'j3�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~Nzq ~Nysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L���uq ~ O   q ~Nq ~
�q ~~w  �sq ~ '�8isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~M=xq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L�ֆouq ~ O   q ~MHw  	sq ~ 'D��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~=�t gainesville:nxq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L�m{Cuq ~ O   q ~=�w  �sq ~ '��7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L�JCOuq ~ O   q ~ Qq ~ �q ~�w  -sq ~ 'w�l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L�"�uq ~ O   q ~"w  �sq ~ 'X^�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L.?��uq ~ O   q ~ Qq ~ �q ~B�w  �sq ~ '��Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L���2uq ~ O   q ~Uw  [sq ~ 'h�Nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ Lx���uq ~ O   q ~ Qq ~ �q ~7w  sq ~ '��{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ft 
arkansas:nxq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L����uq ~ O   q ~fw  Fsq ~ '��usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/�xq ~N�q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~N�sq ~ L��5�uq ~ O   q ~/�q ~ w   isq ~ '�Q6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~O q ~N�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Osq ~ L���uq ~ O   q ~ Qq ~Nq ~ �w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~Oq ~Osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Osq ~ L��Cuq ~ O   q ~$�q ~	�w  zsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/�xq ~Oq ~Osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O sq ~ LZ��Ruq ~ O   q ~/�q ~=w  �sq ~ 'se��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ �t 	madison:nxq ~O'q ~O&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O/sq ~ L1?�uq ~ O   q ~ �w  �sq ~ ' �)[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7@xq ~O6q ~O5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O<sq ~ L���7uq ~ O   q ~7Kt ndw  sq ~ 'z'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	alameda:nxq ~ODq ~OCsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~OLsq ~ L���uq ~ O   q ~�w  gsq ~ '�>�msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~OSq ~ORsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~OYsq ~ L���uq ~ O   q ~ Qq ~ �q ~Fw  3sq ~ 'h�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~]xq ~O`q ~O_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ofsq ~ L�X�uq ~ O   q ~hq ~w  �sq ~ '�zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~8it ewa:nxq ~Omq ~Olsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ousq ~ L �-uq ~ O   q ~8iw  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
richardsont richardson:nxq ~O|q ~O{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O�sq ~ L�^yuq ~ O   q ~O~w  �sq ~ '!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O�sq ~ LB�juq ~ O   q ~�q ~�w  sq ~ ' 8)Csq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~O�sq ~ L 7�uq ~ O   q ~w   0sq ~ '_09sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t san_franciscot san_francisco:nxq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O�sq ~ L"V�uq ~ O   q ~ �q ~		w  �sq ~ '�Jz�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	!xq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~O�sq ~ L i�uq ~ O   q ~ Qq ~w   sq ~ 'I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O�sq ~ L��'uq ~ O   q ~�w  �sq ~ 'r��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~O�sq ~ L\��&uq ~ O   q ~*w   Ysq ~ '�C��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~MHt 	kenosha:nxq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O�sq ~ L�ֆouq ~ O   q ~MHw  �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t tallahassee:nxq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~O�sq ~ L)��uq ~ O   q ~�w  �sq ~ 'M�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#�xq ~O�q ~O�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Psq ~ L���-uq ~ O   q ~ Qq ~#�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~Pq ~Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Psq ~ L<��uq ~ O   q ~Wq ~w  �sq ~ '�BVgsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~><xq ~Pq ~Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Psq ~ LG��Ruq ~ O   q ~*q ~�q ~�w  �sq ~ 'ĕF�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~P"q ~P!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P(sq ~ Ly�)uq ~ O   q ~�q ~ �w  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~P/q ~P.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P5sq ~ L l>uq ~ O   q ~�q ~�w  6sq ~ '��osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-Nxq ~P<q ~P;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~PBsq ~ LFLeuq ~ O   q ~ Qq ~ �q ~-Yw  �sq ~ '��\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~PIq ~PHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~POsq ~ L��ݱuq ~ O   q ~ Qq ~*w  .sq ~ '�_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~PVq ~PUsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P\sq ~ L���uq ~ O   q ~ Qq ~ Rq ~ Sq ~w  �sq ~ 'P7U�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8=xq ~Pcq ~Pbsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Pisq ~ L>��quq ~ O   q ~�w  ysq ~ 's�s9sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Ppq ~Posq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Pvsq ~ L[k�uq ~ O   q ~ Qq ~ �q ~w  	�sq ~ '�7�q ~�sq ~ sq ~ sq ~ J   w   q ~|xq ~P|q ~P{sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~P�sq ~ L^U�uq ~ O   q ~�w  	�sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	phoenix:nxq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ L�}��uq ~ O   q ~�w  	�sq ~ '7b7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ L=�q�uq ~ O   q ~gq ~/q ~0q ~"w  �sq ~ 'Y���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~B�t 	arizona:sxq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ L.���uq ~ O   q ~ Qq ~ Rq ~ Sq ~B�w  	sq ~ '�W�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ L��COuq ~ O   q ~�w   sq ~ '�vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~:xq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ LU���uq ~ O   q ~ Qq ~ �q ~Ew  .sq ~ '��n�q ~$�sq ~ sq ~ sq ~ 
w   q ~�q ~$�xq ~P�q ~P�sq ~ @q ~$�sq ~ G�Uܘ    sq ~ sq ~ J   w   q ~�q ~ �xq ~P�q ~%w   hsq ~ '�|��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ L� ˈuq ~ O   q ~ �q ~�q ~w  ^sq ~ '���rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ L-6�uq ~ O   q ~ Qq ~ �q ~!�q ~!�w  Rsq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~P�sq ~ Lk!�uq ~ O   q ~!�q ~Tw  �sq ~ '6kasq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t ohio:sxq ~P�q ~P�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Qsq ~ L�"�uq ~ O   q ~ Rq ~ Sq ~�w   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~Q
q ~Q	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Qsq ~ L�^Luq ~ O   t americaw  ksq ~ '=)Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~7Kt fargo:nxq ~Qq ~Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q sq ~ L�.}uq ~ O   q ~7Kw  �sq ~ '�)U�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Q'q ~Q&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q-sq ~ L��huq ~ O   q ~ Qq ~ �q ~�q ~�w  sq ~ '��Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~Q4q ~Q3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q:sq ~ L�8l�uq ~ O   q ~-�w  !sq ~ '��� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~QAq ~Q@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~QGsq ~ L����uq ~ O   q ~w  msq ~ '� u�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~QNq ~QMsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~QTsq ~ L�r�uq ~ O   q ~-�q ~Aw  �sq ~ '#hԡsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt springfield_oht springfield_oh:cxq ~Q[q ~QZsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Qdsq ~ L�>2uq ~ O   q ~Fq ~�w  @sq ~ 'h�[\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~Qkq ~Qjsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Qqsq ~ LŊ�uq ~ O   q ~�q ~	bw  �sq ~ '��%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~Qxq ~Qwsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q~sq ~ Lϟkuq ~ O   q ~+Vq ~ Rw  ssq ~ '��`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~&�t 	lincoln:nxq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ L
��=uq ~ O   q ~&�w   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ L�(�uq ~ O   q ~�q ~Uw  sq ~ '�
�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Q�sq ~ L���uq ~ O   t deathw  
sq ~ '�ck�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Q�sq ~ L�b�uq ~ O   q ~w  	�sq ~ '�� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ L 7��uq ~ O   q ~&�w  �sq ~ '����q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~Pq ~ �t 
city:<c,t>xq ~Q�q ~Q�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Q�sq ~ L .��uq ~ O   q ~ �w  	�sq ~ 'a�Z;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ L�>��uq ~ O   q ~�q ~w  �sq ~ ':.s_sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ L�i�uq ~ O   q ~wq ~�q ~�w  	�sq ~ '"HIxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~0t chesapeake:nxq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ LV�vuq ~ O   q ~0w  �sq ~ '�LTsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~Q�q ~Q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Q�sq ~ L7�r�uq ~ O   q ~ Qq ~ �q ~_w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~|xq ~Rq ~R sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Rsq ~ L -��uq ~ O   q ~[w   _sq ~ '��2�q ~�sq ~ sq ~ sq ~ J   w   q ~E�q ~xq ~Rq ~Rsq ~ @q ~�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~Rsq ~ L  �uq ~ O   q ~0�w  
sq ~ '���xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~	�t cambridge:nxq ~Rq ~Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R sq ~ L��Vuq ~ O   q ~	�w  	sq ~ '�G��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	garland:nxq ~R'q ~R&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R/sq ~ L���uq ~ O   q ~�w  �sq ~ '���jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
 xq ~R6q ~R5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R<sq ~ L�x�uq ~ O   q ~ Qq ~ �q ~
q ~
w  �sq ~ 'g�"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~RCq ~RBsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~RIsq ~ L�ʄ�uq ~ O   q ~ �q ~ �q ~"w  0sq ~ '*"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~RPq ~ROsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~RVsq ~ LK�]�uq ~ O   q ~$�q ~	bq ~"w  �sq ~ '暍�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~R]q ~R\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rcsq ~ Ln�(uq ~ O   q ~<q ~ �w  �sq ~ '^�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Rjq ~Risq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Rpsq ~ L�uq ~ O   q ~�q ~ �w  sq ~ '�Vw�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bxq ~Rwq ~Rvsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R}sq ~ L/��uq ~ O   q ~Mq ~�w  �sq ~ ' 0�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~R�sq ~ L 0kOuq ~ O   t givew  	�sq ~ '_ԡ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
dundalk_mdt dundalk_md:cxq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L���uq ~ O   q ~ Qq ~ �q ~&zw  �sq ~ ''=Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L�1�Kuq ~ O   q ~Fw  Wsq ~ 'aVEcsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L--��uq ~ O   q ~ Qq ~ Rq ~ Sq ~"w  sq ~ '#�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L�
uq ~ O   q ~Fq ~w  �sq ~ 'esI�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8|xq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ LsFuq ~ O   q ~8�q ~#Hw  �sq ~ '�02sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8|xq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L�nY�uq ~ O   q ~8�q ~�q ~4w  �sq ~ '�fa�q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~R�q ~R�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~R�sq ~ LRNuq ~ O   q ~7 w  
#sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t nevada:nxq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L�{v�uq ~ O   q ~�w  sq ~ '��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~D�xq ~R�q ~R�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~R�sq ~ L���uq ~ O   q ~D�q ~D�q ~ �w  	nsq ~ '���?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Sq ~Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S
sq ~ L��E�uq ~ O   q ~q ~q ~w  	^sq ~ 'JP��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Sq ~Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ssq ~ L}�Duq ~ O   q ~�q ~�w  (sq ~ '�^isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~Sq ~Ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S$sq ~ Lg�uq ~ O   q ~ Qq ~ Rq ~ Sq ~Mw  �sq ~ '9ca�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/�xq ~S+q ~S*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S1sq ~ L�{�uq ~ O   q ~/�q ~ �w  sq ~ 'Sm�Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+xq ~S8q ~S7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S>sq ~ Lv��uq ~ O   q ~ Qq ~ �q ~ �w  �sq ~ '�?Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~SEq ~SDsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~SKsq ~ L�Ј�uq ~ O   q ~ Qq ~ �q ~!)w  �sq ~ '��d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~SRq ~SQsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~SXsq ~ LQ^4uq ~ O   q ~ �q ~ �w  �sq ~ '*22�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~S_q ~S^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Sesq ~ L�k�uq ~ O   q ~�q ~ �w  �sq ~ 't��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Slq ~Sksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Srsq ~ L�˕�uq ~ O   q ~�q ~�w   �sq ~ '#}q ~�sq ~ sq ~ sq ~ J   w   q ~)xq ~Sxq ~Swsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~S|q ~-�w  	�sq ~ '߃Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ L����uq ~ O   q ~�q ~ Rw   �sq ~ 'W$��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ L\���uq ~ O   q ~�w  sq ~ '��|�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ L.�5uq ~ O   q ~ Qq ~ �q ~Fq ~ �w  3sq ~ 'd�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ L�>�uq ~ O   q ~!�q ~ �w  *sq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7yxq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ LН$�uq ~ O   q ~7�w  Ysq ~ 'Z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ L��1�uq ~ O   q ~ Qq ~ �q ~'w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~S�sq ~ L��]uq ~ O   t smallestw   sq ~ '=���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	yxq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ Ln�"uq ~ O   q ~	�q ~(�w  �sq ~ '�asq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
salton_seat salton_sea:lxq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~S�sq ~ L,�uq ~ O   q ~t saltont seaw  �sq ~ '͞ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~S�q ~S�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L����uq ~ O   q ~q ~=q ~	bw  �sq ~ '�{��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@�xq ~T	q ~Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ LX+�uq ~ O   q ~ Qq ~ �q ~@�w  gsq ~ '.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~F#xq ~Tq ~Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ L��uq ~ O   q ~F.q ~�w  gsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~T#q ~T"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T)sq ~ L�x�uq ~ O   q ~Nq ~�w   �sq ~ '��Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t st_clairt 
st_clair:lxq ~T0q ~T/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T9sq ~ L�|DMuq ~ O   q ~q ~Nq ~w  sq ~ '�6�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'xq ~T@q ~T?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~TFsq ~ L����uq ~ O   q ~ Qq ~ �q ~2w  gsq ~ 'm���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~.t 	georgia:sxq ~TMq ~TLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~TUsq ~ LV"'�uq ~ O   q ~ Qq ~ Rq ~ Sq ~.w  	<sq ~ '�J��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~T\q ~T[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tbsq ~ LS��uq ~ O   q ~ Qq ~ �q ~w  �sq ~ '�e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~Tiq ~Thsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tosq ~ L{�uq ~ O   q ~ Qq ~ �q ~!�w  sq ~ '��+{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"exq ~Tvq ~Tusq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T|sq ~ L��Vuq ~ O   q ~?q ~�w  Vsq ~ '��~sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ L�H	�uq ~ O   q ~[q ~�w  sq ~ '͸��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ LF:�uq ~ O   q ~q ~ww  �sq ~ '  �q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~T�sq ~ L  �uq ~ O   q ~>�w  
 sq ~ '�  �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=�xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ L�m{Cuq ~ O   q ~=�w  ,sq ~ 'A�0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ L�uq ~ O   q ~�q ~ �w  �sq ~ '`3�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t san_joset 
san_jose:nxq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ L g�Wuq ~ O   q ~ �q ~Nw  ;sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ LJ�buq ~ O   q ~ Qq ~
q ~ �w  Ssq ~ '��G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~P�xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ L�Ų>uq ~ O   q ~B�w  ysq ~ '�ƈ>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@�xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ L�:�Wuq ~ O   q ~q ~#w  �sq ~ '��Asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~T�q ~T�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~T�sq ~ Lɐ�'uq ~ O   q ~ Rq ~ Sq ~
�q ~
�w   �sq ~ '��Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Uq ~Usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U	sq ~ L�f�Suq ~ O   q ~ Qq ~ �q ~%w  �sq ~ 'o��Osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4xq ~Uq ~Usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Usq ~ Lװ/�uq ~ O   q ~ Qq ~ �q ~?w  �sq ~ ' 3~�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Uq ~1w  	�sq ~ '�Rxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~7t koolaupoko:nxq ~U#q ~U"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U+sq ~ LlMG�uq ~ O   q ~7w  �sq ~ '�
��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3�xq ~U2q ~U1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U8sq ~ L����uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '<H��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
brockton:nxq ~U?q ~U>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~UGsq ~ L��juq ~ O   q ~�w  �sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t east_los_angelest east_los_angeles:nxq ~UNq ~UMsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~UWsq ~ L~�Zuq ~ O   q ~gq ~/q ~0w   �sq ~ '�*UHq ~�sq ~ sq ~ sq ~ J   w   q ~Hxq ~U]q ~U\sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~Uasq ~ L�8�euq ~ O   t heightw  
sq ~ 'v��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9�xq ~Uiq ~Uhsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Uosq ~ LmyRXuq ~ O   q ~
�q ~9�q ~"w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ht birmingham:nxq ~Uvq ~Uusq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U~sq ~ L��b�uq ~ O   q ~Hw  >sq ~ '>�v�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/4xq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ Lʌ'�uq ~ O   q ~ Qq ~ Rq ~ Sq ~
�q ~�w  {sq ~ 'S�(�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L[5�uq ~ O   q ~ Qq ~ Rq ~ Sq ~w  (sq ~ '�A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6�xq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L"tK;uq ~ O   q ~6�q ~ �w  Ssq ~ '�"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t montgomery:nxq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L���uq ~ O   q ~�w  Isq ~ '���Zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*xq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L0���uq ~ O   q ~ Qq ~ �q ~ q ~5w  �sq ~ 'x��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L���uq ~ O   q ~4q ~+w  �sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t west_covinat west_covina:nxq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L���#uq ~ O   q ~q ~=w  :sq ~ 'q�:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ LU�uq ~ O   q ~�q ~w  Isq ~ '�Z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~*t carson:nxq ~U�q ~U�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~U�sq ~ L�|=|uq ~ O   q ~*w   �sq ~ 'P/�q ~�sq ~ sq ~ sq ~ J   w   q ~;xq ~V q ~U�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Vsq ~ L�mlIuq ~ O   t capitalsw  	�sq ~ '7qG�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<jxq ~Vq ~Vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Vsq ~ L�Q��uq ~ O   q ~"Nq ~5w  	[sq ~ '���!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Vq ~Vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Vsq ~ L\ڤuq ~ O   q ~�w  �sq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~3t minnesota:nxq ~V&q ~V%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V.sq ~ L8�quq ~ O   q ~3w  �sq ~ 'Ĭ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~V5q ~V4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V;sq ~ L�;��uq ~ O   q ~�q ~�t nvw  �sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t hollywood:nxq ~VCq ~VBsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~VKsq ~ LV��}uq ~ O   q ~�w  dsq ~ 'i��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~"	t 	bayonne:nxq ~VRq ~VQsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~VZsq ~ L��.uq ~ O   q ~"	w  asq ~ '>��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)4xq ~Vaq ~V`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Vgsq ~ Lw2�uq ~ O   q ~)?w  	�sq ~ '�D�zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	!xq ~Vnq ~Vmsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~Vtsq ~ L c��uq ~ O   q ~q ~3w   :sq ~ '&F��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~V{q ~Vzsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ L�a2�uq ~ O   q ~2�q ~�q ~�w  �sq ~ '���;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t rhode_island:nxq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ L�)��uq ~ O   q ~�q ~�w  �sq ~ 'U��Wq ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~V�q ~V�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~V�sq ~ L�-v]uq ~ O   t containsw  
sq ~ '�~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ L���iuq ~ O   q ~ Qq ~ �q ~�q ~�w  �sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ LayԲuq ~ O   q ~�q ~�q ~ w  �sq ~ 'Ӵ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~7it 	modesto:nxq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ LI!��uq ~ O   q ~7iw  |sq ~ '1�@�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ L5�nquq ~ O   q ~ Qq ~ �q ~�w  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*$xq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ L����uq ~ O   q ~�t idw  wsq ~ '�+�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~V�sq ~ L���uq ~ O   q ~�w  
Rsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~V�q ~V�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~V�sq ~ Le�j�uq ~ O   q ~Fw  �sq ~ '("q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~V�sq ~ L(��uq ~ O   t populousw  	�sq ~ 'lN��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Wq ~Wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W
sq ~ L���uq ~ O   q ~w  �sq ~ 'U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Wq ~Wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Wsq ~ L���uq ~ O   q ~�w  �sq ~ '�ֳ+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~Wq ~Wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W$sq ~ L��;uq ~ O   q ~wq ~�w  Osq ~ '�	Fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~W+q ~W*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W1sq ~ L�"U�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�[z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~W8q ~W7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W>sq ~ LG�quq ~ O   q ~ Rq ~ Sq ~�w  #sq ~ '?��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~WEq ~WDsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~WKsq ~ L�%Muq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  �sq ~ '�9#q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0sq ~ �?���t 	<e,<n,t>>q ~ <sq ~ ��6�t <n,t>q ~�q ~ �t namedt named:<e,<n,t>>xq ~WQq ~WPsq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~W\sq ~ L;׆uq ~ O   t namesw  
;sq ~ '�c� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Wdq ~Wcsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Wjsq ~ L:KMuq ~ O   q ~�w  �sq ~ '�\nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Wqq ~Wpsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Wwsq ~ L�5huq ~ O   q ~ �q ~�w  	bsq ~ '�W'bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~W~q ~W}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L�7Ouq ~ O   q ~B�w  �sq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt 
mount_sillt mount_sill:mxq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L��)=uq ~ O   q ~ zt sillw  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L��yuq ~ O   q ~�q ~�w  �sq ~ ')���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ LHR{cuq ~ O   q ~ Qq ~�q ~�w  Msq ~ '�R�9sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,{xq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L�Q��uq ~ O   q ~ Qq ~ �q ~'0w  tsq ~ 'Y^:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L�"�uq ~ O   q ~ Qq ~ �q ~�w  Ssq ~ '�pA�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Uxq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L��,�uq ~ O   q ~ �q ~`q ~ �w  5sq ~ '^] �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"sxq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L����uq ~ O   q ~�q ~Aw  Wsq ~ 'k��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Exq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~W�sq ~ L��uq ~ O   q ~Dw   .sq ~ '��Bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~exq ~W�q ~W�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~W�sq ~ L�Z�uq ~ O   q ~pq ~Uq ~�w  jsq ~ '��C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
santa_rosat santa_rosa:nxq ~Xq ~Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Xsq ~ L��|~uq ~ O   q ~ q ~w   �sq ~ 'vU&Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ t 
virginia:nxq ~Xq ~Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Xsq ~ L\�Mcuq ~ O   q ~ w  {sq ~ '�Y�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~M_xq ~X#q ~X"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X)sq ~ Lm��uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '[y�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'t durham:nxq ~X0q ~X/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X8sq ~ L�J�1uq ~ O   q ~'w  �sq ~ '���Fq ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~X>q ~X=sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~XBsq ~ L��auq ~ O   q ~Ww  
Vsq ~ '_U@�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Rxq ~XIq ~XHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~XOsq ~ LŅ��uq ~ O   q ~]q ~	q ~ gw  �sq ~ ')��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~XVq ~XUsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X\sq ~ L 2�Kuq ~ O   q ~1w  �sq ~ 'r��@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~Xcq ~Xbsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Xisq ~ L��-]uq ~ O   q ~B�q ~iw  �sq ~ '|��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~Xpq ~Xosq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Xvsq ~ L���uq ~ O   q ~ Rq ~ Sq ~�q ~�w  ]sq ~ ' �q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~X~sq ~ L y�uq ~ O   t allw  	�sq ~ '&��\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~wxq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L���>uq ~ O   q ~�q ~�q ~�q ~�w  sq ~ '�ѧ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+rxq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L�+��uq ~ O   q ~+}q ~�w  	sq ~ '���;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L���uq ~ O   q ~�q ~w   �sq ~ '�'��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L`�r�uq ~ O   q ~�q ~�w  �sq ~ '���[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t thousand_oakst thousand_oaks:nxq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L �{|uq ~ O   q ~D�q ~D�w   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ Lir�Auq ~ O   q ~ Rq ~ Sq ~#w  	�sq ~ '�<��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8Mxq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ Lr�+uq ~ O   q ~ Qq ~8Xq ~ �w  	Psq ~ '`:��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'�t 	meriden:nxq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L8�huq ~ O   q ~'�w  &sq ~ '�7rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~K�xq ~X�q ~X�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~X�sq ~ L�pHuq ~ O   q ~ Rq ~ Sq ~�w  �sq ~ '�=q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~Ysq ~ L���uq ~ O   q ~ Rw  	�sq ~ 'Cr88sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Yq ~Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~Ysq ~ L���uq ~ O   q ~ Rw   `sq ~ '�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~Yq ~Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ysq ~ L�|�fuq ~ O   q ~Fw  �sq ~ '<���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~wxq ~Y"q ~Y!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y(sq ~ L]�uq ~ O   q ~�w  	xsq ~ 'p���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"exq ~Y/q ~Y.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y5sq ~ L��u�uq ~ O   q ~ Qq ~ �q ~?w  �sq ~ '7/�)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~Y<q ~Y;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~YBsq ~ Lk�c�uq ~ O   q ~�w  bsq ~ '�rrsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~YIq ~YHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~YOsq ~ Lo�uq ~ O   q ~ Rq ~ Sq ~"w  �sq ~ '
{��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~YVq ~YUsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y\sq ~ L�}��uq ~ O   q ~�w  �sq ~ '�_`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1�xq ~Ycq ~Ybsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Yisq ~ Lo�uq ~ O   q ~ �q ~1�q ~ �w  sq ~ '�6Dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Ypq ~Yosq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Yvsq ~ L�"3uq ~ O   q ~ Qq ~ �q ~�w   �sq ~ '�,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~,t 	vallejo:nxq ~Y}q ~Y|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L��]uq ~ O   q ~,w  �sq ~ '�وsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L��?^uq ~ O   q ~�q ~�w   �sq ~ '�5w�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L�d�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�l��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t jersey_cityt jersey_city:nxq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L�X��uq ~ O   q ~Fq ~ �w  rsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~4t macon:nxq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L-��uq ~ O   q ~4w  sq ~ 'aD�q ~�sq ~ sq ~ sq ~ J   w   q ~xq ~Y�q ~Y�sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L ��uq ~ O   q ~"w  
@sq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~"t 	florida:nxq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L�X�uq ~ O   q ~"w  �sq ~ '~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#yxq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ LC�guq ~ O   q ~�q ~#�q ~�w  Bsq ~ 'd�ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L���uq ~ O   q ~Uq ~
�q ~ Rw  sq ~ '�,�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
 xq ~Y�q ~Y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Y�sq ~ L]�uq ~ O   q ~
q ~
q ~ �w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~8�t manchester:nxq ~Zq ~Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Zsq ~ L :�uq ~ O   q ~8�w  �sq ~ '�G}8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Et 
paterson:nxq ~Zq ~Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Zsq ~ LIw@uq ~ O   q ~Ew  �sq ~ 'Rmu8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Z#q ~Z"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z)sq ~ L���uq ~ O   q ~�w  sq ~ '�؆�q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~Z/q ~Z.sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~Z3sq ~ LĤtuq ~ O   t 	borderingw  	�sq ~ '�s+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~K�xq ~Z;q ~Z:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ZAsq ~ L��uq ~ O   q ~�q ~ Rw  Zsq ~ '�zX�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
fall_rivert fall_river:nxq ~ZHq ~ZGsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ZQsq ~ LC�uq ~ O   q ~	Pq ~ �w   vsq ~ 'g�>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~ZXq ~ZWsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z^sq ~ LZh�,uq ~ O   q ~ Qq ~ �q ~�w  sq ~ '憟�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~Zeq ~Zdsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Zksq ~ Lp`uq ~ O   q ~!�q ~"w  �sq ~ 'gw��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~MNxq ~Zrq ~Zqsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Zxsq ~ L,|uq ~ O   q ~ Qq ~MYq ~ �w  Wsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9�xq ~Zq ~Z~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�Q[�uq ~ O   q ~ �q ~9�q ~"w  zsq ~ '|�qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4xq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�g~iuq ~ O   q ~?q ~.w  	|sq ~ 'W���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�uq ~ O   q ~ Qq ~ �q ~ww  �sq ~ '��4xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~B�t 	arizona:nxq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�Ų>uq ~ O   q ~B�w  9sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t kansas:nxq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�!/Kuq ~ O   q ~w  1sq ~ '5�;Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"-xq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L£L)uq ~ O   q ~{q ~�w  [sq ~ 'P��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�I�uq ~ O   q ~�q ~ �w  Lsq ~ '$���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ Lag��uq ~ O   q ~ Qq ~ Rq ~ Sq ~ �w  �sq ~ '��j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Z�sq ~ L�t�guq ~ O   q ~ Qq ~�q ~�q ~ �w  sq ~ 'V^�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt springfield_sdt springfield_sd:cxq ~Z�q ~Z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[sq ~ L���uq ~ O   q ~Fq ~
�q ~
�w  �sq ~ '�*$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~[q ~[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[sq ~ L�aWAuq ~ O   q ~!�q ~!�w  'sq ~ '�PR2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~[q ~[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[sq ~ L��Izuq ~ O   q ~ Rq ~ Sq ~Sw  �sq ~ 'Z:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~["q ~[!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[(sq ~ L�B�buq ~ O   q ~�q ~�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~(.t 	yonkers:nxq ~[/q ~[.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[7sq ~ L�|5quq ~ O   q ~(.w  sq ~ '��psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~->xq ~[>q ~[=sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[Dsq ~ L�8��uq ~ O   q ~�w  rsq ~ '��� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt omaha_net 
omaha_ne:cxq ~[Kq ~[Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[Tsq ~ L�� uq ~ O   q ~ Qq ~ �t omahaw  sq ~ 'S�1�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~R�xq ~[\q ~[[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[bsq ~ Lw�.wuq ~ O   q ~&zw  Dsq ~ '�i�(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*Pxq ~[iq ~[hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[osq ~ L��uq ~ O   q ~*[q ~*\w  dsq ~ '��ߘsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6#xq ~[vq ~[usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[|sq ~ LK0uq ~ O   q ~�q ~�q ~Tw  )sq ~ 'ej��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Irxq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ L��H�uq ~ O   q ~I}q ~ gw  �sq ~ 'm�o5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7^xq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ L�?�Muq ~ O   q ~7iq ~"w  �sq ~ 'V��q ~�sq ~ sq ~ sq ~ 
w   q ~	!q ~1vxq ~[�q ~[�sq ~ @q ~�sq ~ G���    sq ~ sq ~ J   w   q ~	,q ~ <xq ~[�q ~�w   esq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ L�b�uq ~ O   q ~ Qq ~ �q ~ �q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ Lㆺuq ~ O   q ~ Qq ~ �q ~w  �sq ~ '�R�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt richmond_vat richmond_va:cxq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ L��FXuq ~ O   q ~ Qq ~ �q ~qw  �sq ~ 'g_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ LO2�]uq ~ O   q ~w  Gsq ~ '�X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ L*���uq ~ O   q ~"q ~ Rw   �sq ~ '�W�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
$xq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ L��/uq ~ O   q ~
/q ~ �w  8sq ~ ',��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~#t 
colorado:nxq ~[�q ~[�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~[�sq ~ Lڄ�uq ~ O   q ~#w  Vsq ~ '�ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~TNxq ~\q ~\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\sq ~ L�L�uq ~ O   q ~.w  �sq ~ '��][sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~\q ~\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\sq ~ L�<�uq ~ O   q ~ Qq ~ �q ~	�w  ;sq ~ '�z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*$xq ~\q ~\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\%sq ~ L�*�uq ~ O   q ~�q ~gw  �sq ~ '�E;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~\,q ~\+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\2sq ~ L��6 uq ~ O   q ~Xw  ~sq ~ '�Ħ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~\9q ~\8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\?sq ~ L��]uq ~ O   q ~,w  xsq ~ '�-7q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~\Gsq ~ L���uq ~ O   t 	populatedw  	�sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
livonia_mit livonia_mi:cxq ~\Oq ~\Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\Xsq ~ LU�,uq ~ O   q ~=Oq ~Tw  )sq ~ '��w8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8-xq ~\_q ~\^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\esq ~ LVm�uq ~ O   q ~�q ~�q ~"w  5sq ~ '�^��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~\lq ~\ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\rsq ~ L�uq ~ O   q ~Nq ~Ow  sq ~ '��j/sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt portland_met portland_me:cxq ~\yq ~\xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ LIX�@uq ~ O   q ~_q ~ >w  �sq ~ '���usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~?axq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ L���Quq ~ O   q ~8�q ~5w  =sq ~ 'ƋOmsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A@xq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ L?<�]uq ~ O   q ~AKq ~�w  sq ~ '��Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_south_buttresst mount_south_buttress:mxq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ LҜ�uq ~ O   q ~ zq ~
�t buttressw  �sq ~ '3'@]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8^xq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ L�61�uq ~ O   q ~8iq ~w  �sq ~ 'Y���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ L�uq ~ O   q ~_q ~�w  �sq ~ '/�-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ Ls<�Luq ~ O   q ~q ~�w  Ksq ~ '��U8q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~\�q ~\�sq ~ @q ~ �sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�q ~ �w   [sq ~ 'A9��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ L��tuq ~ O   q ~Cw  Jsq ~ '��|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt kettering_oht kettering_oh:cxq ~\�q ~\�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~\�sq ~ Lĳ;�uq ~ O   q ~ Qq ~ �t 	ketteringw  1sq ~ ';��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~&t waterford:nxq ~]q ~] sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]	sq ~ L�Dn�uq ~ O   q ~&w  �sq ~ '�}8.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~]q ~]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~]sq ~ L��5�uq ~ O   t lowestw   Csq ~ '=���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$6xq ~]q ~]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]$sq ~ Li��uq ~ O   q ~ Qq ~$Aw  �sq ~ '�.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[�xq ~]+q ~]*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]1sq ~ L����uq ~ O   q ~qw  Esq ~ '_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~]8q ~]7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]>sq ~ L� �puq ~ O   q ~ Qq ~�q ~�w  �sq ~ '��`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~]Eq ~]Dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]Ksq ~ L@e��uq ~ O   q ~!�w  psq ~ '��1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/yxq ~]Rq ~]Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]Xsq ~ L����uq ~ O   q ~ Qq ~ �q ~/�w  5sq ~ 'u���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'Pxq ~]_q ~]^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]esq ~ L��uq ~ O   q ~'[q ~w  �sq ~ '�m��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~]lq ~]ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]rsq ~ LEK4uq ~ O   q ~"q ~ Rw   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
warwick_rit warwick_ri:cxq ~]yq ~]xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ L)�O�uq ~ O   q ~q ~�q ~�w  �sq ~ 'h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ L����uq ~ O   q ~�q ~ �w  �sq ~ '\o�asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8=xq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ LK D�uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '���q ~	sq ~ sq ~ sq ~ 
w   q ~�q ~	!xq ~]�q ~]�sq ~ @q ~	'sq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~]�q ~	.w   Nsq ~ 'kÛsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[Lxq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ L×��uq ~ O   q ~[Wq ~,�w  �sq ~ 'r1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t terre_hautet terre_haute:nxq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ LўfYuq ~ O   q ~�q ~�w  7sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
mille_lacst mille_lacs:lxq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ L~Iuq ~ O   q ~t millet lacsw  �sq ~ 'u�$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ L��Z�uq ~ O   q ~ Qq ~ �q ~Dw  	sq ~ '�}`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Ixq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ Lx7ȧuq ~ O   q ~1�q ~w  �sq ~ 'ٚ)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~/�t 	norfolk:nxq ~]�q ~]�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~]�sq ~ L~��uq ~ O   q ~/�w  �sq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~_xq ~^q ~^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^	sq ~ Lbj�uq ~ O   q ~jq ~5w  sq ~ ' �Tq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~^sq ~ L zuq ~ O   t andw  
Asq ~ '�F��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~^q ~^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^sq ~ L��FXuq ~ O   q ~ Qq ~ �q ~qw  asq ~ '��?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~^&q ~^%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^,sq ~ L�.��uq ~ O   q ~ Qq ~ �q ~ �q ~ �w  	�sq ~ 'v-�qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~^3q ~^2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^9sq ~ L�*#9uq ~ O   q ~�w  �sq ~ 'u˒�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t plano:nxq ~^@q ~^?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^Hsq ~ L\ڤuq ~ O   q ~�w  �sq ~ 'G5�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+xq ~^Oq ~^Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^Usq ~ L>-yuq ~ O   q ~ �w  �sq ~ ' 1�Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~^\q ~^[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~^bsq ~ L 1�	uq ~ O   q ~t feetw   &sq ~ '�W�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~^jq ~^isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^psq ~ L�l�uq ~ O   q ~fq ~Tw  �sq ~ 'y^�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt sioux_falls_sdt sioux_falls_sd:cxq ~^wq ~^vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ L0��uq ~ O   q ~Uq ~Et sdw   �sq ~ '�	N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~\�t kettering:nxq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ L�z�9uq ~ O   q ~\�w  Fsq ~ '��f;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ L���uq ~ O   q ~�q ~=w  �sq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t eugene:nxq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ L���uq ~ O   q ~�w  �sq ~ '~��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ L+u*uq ~ O   q ~_w  �sq ~ '7umVsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\xq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ LG��Yuq ~ O   q ~ Qq ~ �q ~/q ~0w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3xq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ LH���uq ~ O   q ~~q ~�w  Lsq ~ '��q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t yellowstone_rivert yellowstone_river:rxq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ Lp O�uq ~ O   t yellowstoneq ~ �w  sq ~ '�&��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~D�xq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ L�#�uq ~ O   q ~D�q ~D�q ~"w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"=xq ~^�q ~^�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~^�sq ~ Lc��uq ~ O   q ~�q ~"w  gsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%	xq ~_q ~_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_sq ~ LPZ��uq ~ O   q ~%q ~ gw  �sq ~ '��;	q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~_q ~_sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~_sq ~ L�;$uq ~ O   t lengthw  
sq ~ ' �C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~_q ~_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_#sq ~ Li<#�uq ~ O   q ~ �q ~�q ~#w  �sq ~ '|�,�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\�xq ~_*q ~_)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_0sq ~ LVަuq ~ O   q ~\�q ~	�w  	5sq ~ 'J��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)4xq ~_7q ~_6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_=sq ~ L�j|Auq ~ O   q ~ Qq ~ �q ~)?w  �sq ~ '1��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~+t utica:nxq ~_Dq ~_Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_Lsq ~ L��uq ~ O   q ~+w  msq ~ '�Ovsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~_Sq ~_Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_Ysq ~ L 6`-uq ~ O   q ~ Qq ~hw  <sq ~ '�*��q ~sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~__q ~_^sq ~ @q ~sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~_cq ~w   sq ~ '3�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~G�xq ~_hq ~_gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_nsq ~ LU�W�uq ~ O   q ~�w  �sq ~ '�'usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~_uq ~_tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_{sq ~ L
Kt�uq ~ O   q ~�q ~"w  isq ~ 'U]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L���luq ~ O   q ~ Qq ~ �q ~[w  sq ~ 'H�.^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~wxq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ LiU\suq ~ O   q ~ Qq ~ �q ~�w  *sq ~ '�ޤ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
oklahoma:nxq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L�x�uq ~ O   q ~�w  usq ~ 'T�.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6#xq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L� ߥuq ~ O   q ~ Qq ~ �q ~�q ~�w  Tsq ~ '����q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~_�sq ~ L��.�uq ~ O   q ~Iw  
sq ~ 'azT<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L 8
 uq ~ O   q ~ Qq ~"w  �sq ~ '
}��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L���uq ~ O   q ~ Qq ~ �q ~Xw  bsq ~ '�,J(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Rxq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L)\�/uq ~ O   q ~]q ~	q ~Tw  �sq ~ ''��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ Lh�-�uq ~ O   q ~�q ~�q ~�w  	{sq ~ 'c�s|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~_�q ~_�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~_�sq ~ L�NB�uq ~ O   q ~ Qq ~ �w  �sq ~ 'y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6xq ~`q ~` sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`sq ~ L��i`uq ~ O   q ~ Qq ~ �q ~
/w  �sq ~ 'l/�?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~`q ~`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`sq ~ L��.�uq ~ O   q ~ Qq ~ �q ~#w  �sq ~ '�>͜sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t truet true:txq ~`q ~`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  T    sq ~ sq ~ J   w   q ~ �xq ~`$sq ~ L�Jpuq ~ O   t areq ~1%w   bsq ~ 'g4�Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~`,q ~`+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`2sq ~ LNЛWuq ~ O   q ~�q ~ w  Ysq ~ '�6Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~jxq ~`9q ~`8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`?sq ~ L��uq ~ O   q ~ Qq ~ �q ~uw  {sq ~ '��/�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Hxq ~`Fq ~`Esq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`Lsq ~ Lk�C�uq ~ O   q ~Sw   �sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~`Sq ~`Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`Ysq ~ L�}�uq ~ O   q ~�q ~w  sq ~ '��1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~``q ~`_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`fsq ~ LGz\1uq ~ O   q ~q ~
q ~w  ~sq ~ 'j��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~`mq ~`lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`ssq ~ L �Wuq ~ O   q ~2�q ~�q ~�w  vsq ~ '�)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\zxq ~`zq ~`ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L7�r�uq ~ O   q ~ Qq ~ �q ~_w  �sq ~ '�狽sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L�I�uq ~ O   q ~�w  �sq ~ '^[�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~R�xq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L���^uq ~ O   q ~&zq ~&cw  �sq ~ 'դ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L�`��uq ~ O   q ~�q ~ gw  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Yxq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ LŮ�uq ~ O   q ~ fw  	sq ~ '�v�<q ~�sq ~ sq ~ sq ~ J   w   q ~WRxq ~`�q ~`�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~`�sq ~ L�yg�uq ~ O   t calledw  	�sq ~ '��.	sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-Nxq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L:��uq ~ O   q ~-Yw  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~18xq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L��^9uq ~ O   q ~1Cq ~Uq ~�w  �sq ~ '��.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L�]�uq ~ O   q ~ Qq ~ �q ~$�w  rsq ~ 'vv4�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)�xq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~`�sq ~ L�~~uq ~ O   q ~ Qq ~ �q ~ w  �sq ~ 'z���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t fort_lauderdalet fort_lauderdale:nxq ~`�q ~`�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~asq ~ Lb�uq ~ O   q ~ �q ~9�w  �sq ~ '�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~a
q ~a	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~asq ~ L�{v�uq ~ O   q ~�w  �sq ~ '���q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~asq ~ L��tjuq ~ O   q ~$Ow  
"sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~aq ~asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a%sq ~ L��eEuq ~ O   q ~�q ~ Rw  �sq ~ '�]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t newport_newst newport_news:nxq ~a,q ~a+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a5sq ~ LS9`�uq ~ O   q ~3q ~'�w  sq ~ '�;1Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t mississippi:nxq ~a<q ~a;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~aDsq ~ LY�!+uq ~ O   q ~�w  sq ~ '"T$ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Hxq ~aKq ~aJsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~aQsq ~ L�B8�uq ~ O   q ~Sq ~ gw  �sq ~ '�I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~wxq ~aXq ~aWsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a^sq ~ LJ�uq ~ O   q ~�q ~�q ~ �w  �sq ~ 'd�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~}t 
nebraska:sxq ~aeq ~adsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~amsq ~ L/E�uq ~ O   q ~}w  �sq ~ '
�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~%\t boston:nxq ~atq ~assq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a|sq ~ L��&uq ~ O   q ~%\w  _sq ~ '3u��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L�jO�uq ~ O   q ~ Qq ~ �q ~Fw  �sq ~ '�߯�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t lafayette:nxq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L�KL�uq ~ O   q ~�w  �sq ~ 'L�S|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L���uq ~ O   q ~#q ~B�w  2sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L�u��uq ~ O   q ~�w  Vsq ~ '�c�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L�@z�uq ~ O   q ~ �q ~�q ~"w  �sq ~ '-4{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ Lxouq ~ O   q ~'q ~_w  sq ~ '�Ɇ8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ Lv�uq ~ O   q ~Nq ~Oq ~�w   ~sq ~ '��_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~nxq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L��h�uq ~ O   q ~ Qq ~ �q ~yw  �sq ~ 'w�Yxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~"t california:nxq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~a�sq ~ L�"�uq ~ O   q ~"w  +sq ~ '48Ըsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~a�q ~a�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bsq ~ Lb]_ruq ~ O   q ~&�q ~�q ~(�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
south_gatet south_gate:nxq ~b	q ~bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bsq ~ L���~uq ~ O   q ~
�q ~9�w  5sq ~ '�[|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"-xq ~bq ~bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bsq ~ L~�lXuq ~ O   q ~{w  �sq ~ '�uW�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~b&q ~b%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b,sq ~ L��+uq ~ O   q ~q ~ �w  �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~A-t 	anaheim:nxq ~b3q ~b2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b;sq ~ L�y>�uq ~ O   q ~A-w  Jsq ~ 'k��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~bBq ~bAsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bHsq ~ Lg�zuq ~ O   q ~Tw  �sq ~ '�P�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~bOq ~bNsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bUsq ~ LL�?0uq ~ O   q ~ Qq ~ �q ~!�w  	�sq ~ '܎!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	yxq ~b\q ~b[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~bbsq ~ L+�uq ~ O   q ~	�q ~�q ~Fw  �sq ~ '5IA<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t powder_rivert powder_river:rxq ~biq ~bhsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~brsq ~ LŨ�Huq ~ O   q ~ Qt powderw  �sq ~ 'n$��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~bzq ~bysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L�[��uq ~ O   q ~!�q ~!�q ~ �w  �sq ~ '�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L���euq ~ O   q ~ Qq ~ Rq ~ Sq ~�q ~Fw   �sq ~ 'w�h q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~b�q ~b�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~b�sq ~ L  &uq ~ O   t gow  
6sq ~ 'b���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ Lv�K�uq ~ O   q ~Nq ~q ~�w  �sq ~ '� e<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#hxq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L��5uq ~ O   q ~ Qq ~#sq ~ �w  Qsq ~ 'HM�q ~�sq ~ sq ~ sq ~ J   w   q ~Axq ~b�q ~b�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~b�q ~+$w  	�sq ~ '1K��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ Lk�Quq ~ O   q ~�q ~	�w  �sq ~ ' dB�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L��uq ~ O   q ~Wq ~ �w  �sq ~ '}Q8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	fremont:nxq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L���uq ~ O   q ~�w  Rsq ~ 'P�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~^t fayetteville:nxq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L.���uq ~ O   q ~^w  Msq ~ '	T��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~b�q ~b�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~b�sq ~ L�N-xuq ~ O   q ~�q ~�w  �sq ~ ' �88sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t worcester:nxq ~cq ~csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~csq ~ L3���uq ~ O   q ~�w  �sq ~ '<Ҧsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~cq ~csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~csq ~ Ln��`uq ~ O   q ~�w  >sq ~ ']�ppsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t niobrara_rivert niobrara_river:rxq ~c"q ~c!sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c+sq ~ L�Q��uq ~ O   q ~ Qt niobraraq ~ �w  �sq ~ '�b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~c3q ~c2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c9sq ~ L5-�uq ~ O   q ~�w  �sq ~ '�suPsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'axq ~c@q ~c?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~cFsq ~ L��GKuq ~ O   q ~'lq ~ �w  	�sq ~ '�W��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~jxq ~cMq ~cLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~cSsq ~ L�E�uq ~ O   q ~uw  Nsq ~ '՘sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~6�t riverside:nxq ~cZq ~cYsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~cbsq ~ L���uq ~ O   q ~6�w   sq ~ 'Bh�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~[Wt omaha:nxq ~ciq ~chsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~cqsq ~ LO6�uq ~ O   q ~[Ww  gsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'lt 	lubbock:nxq ~cxq ~cwsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L[9,uq ~ O   q ~'lw  	qsq ~ '`X��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ LN�H&uq ~ O   q ~ Qq ~ �q ~2�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ Lˁ�auq ~ O   q ~�w  sq ~ 'R��|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L��'uq ~ O   q ~ Qq ~'�w  �sq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~0�t nashville:nxq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L�N�Huq ~ O   q ~0�w  sq ~ '�.��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0xq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L�	�uq ~ O   q ~ q ~;q ~"w  �sq ~ '�抉q ~�sq ~ sq ~ sq ~ J   w   q ~Zxq ~c�q ~c�sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L���@uq ~ O   q ~!�w  	�sq ~ '���\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^xxq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ LZ�o�uq ~ O   q ~Uq ~Eq ~
�q ~
�w  �sq ~ '	Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~<�t toledo:nxq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L�@��uq ~ O   q ~<�w  �sq ~ '�UMsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~c�sq ~ L�lֹuq ~ O   q ~aq ~�w  	%sq ~ ' ʘ[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~c�q ~c�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ L#C-uq ~ O   q ~+�q ~�w  sq ~ 'H�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t overland_parkt overland_park:nxq ~d
q ~d	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ L�(��uq ~ O   q ~oq ~pw  	ssq ~ '�A"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t st_francis_rivert st_francis_river:rxq ~dq ~dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d#sq ~ L��r�uq ~ O   q ~Nt francisq ~ �w  sq ~ '�NI�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~d,sq ~ L�M�suq ~ O   q ~�w  
Zsq ~ '�
'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~d3q ~d2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d9sq ~ LŢ��uq ~ O   q ~qq ~pw  	�sq ~ '�i�q ~�sq ~ sq ~ sq ~ J   w   q ~�q ~ �xq ~d?q ~d>sq ~ @q ~�sq ~ G�Uܘ    sq ~ sq ~ J   w   q ~�q ~ �xq ~dCsq ~ L  �uq ~ O   q ~>�w  
Lsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/	xq ~dJq ~dIsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dPsq ~ L�Ͻ�uq ~ O   q ~/q ~ gw  !sq ~ 'XbL�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~dWq ~dVsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d]sq ~ Lk�C�uq ~ O   q ~Sw  �sq ~ 'PJ�}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~ddq ~dcsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~djsq ~ L��.uq ~ O   q ~"	w  �sq ~ 'Ԛ �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8q ~�t massachusetts:sxq ~dqq ~dpsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dysq ~ LLwHvuq ~ O   q ~ Rq ~ Sq ~�w  �sq ~ '�Dt�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~d�q ~dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ LgB,iuq ~ O   q ~�q ~Eq ~w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L*S�suq ~ O   q ~�q ~ �w  sq ~ '#4ٻsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Q\xq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L�
Luq ~ O   q ~Fq ~	�w  �sq ~ '��M�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L���uq ~ O   q ~�q ~�q ~ �w   rsq ~ '!w�Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>�xq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L��uq ~ O   q ~�w  ?sq ~ '�Xc�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~]zxq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L/ �uq ~ O   q ~q ~�w  Dsq ~ '�'8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t albuquerque:nxq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L��luq ~ O   q ~�w  ?sq ~ ' q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~d�sq ~ L ��uq ~ O   q ~w  	�sq ~ '�l�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~~xq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ L�BVjuq ~ O   q ~�q ~�q ~w  �sq ~ '�3)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~]zxq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~d�sq ~ LC	��uq ~ O   q ~w   sq ~ 'YՎCsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~d�q ~d�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~esq ~ L����uq ~ O   q ~ Qq ~ Rq ~ Sq ~w  Zsq ~ 'a-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Mxq ~eq ~esq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~esq ~ L��5uq ~ O   q ~ Qq ~ �q ~Xw  �sq ~ '	��2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~eq ~esq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~esq ~ Lbj&uq ~ O   q ~ Qq ~ �q ~w  �sq ~ '�L��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[Lxq ~e&q ~e%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e,sq ~ L��~�uq ~ O   q ~[Wq ~}w  �sq ~ 'ˈz�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t provo:nxq ~e3q ~e2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e;sq ~ L_�duq ~ O   q ~�w  �sq ~ 'K�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_harvardt mount_harvard:mxq ~eBq ~eAsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~eKsq ~ L��uq ~ O   q ~ zt harvardw  �sq ~ '�C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~eSq ~eRsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~eYsq ~ Lׄ�{uq ~ O   q ~ Qq ~�q ~ �w  fsq ~ 'p˰�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_torreyst mount_torreys:mxq ~e`q ~e_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~eisq ~ L|��Kuq ~ O   q ~ zt torreysw  sq ~ 'C�Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6#xq ~eqq ~epsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ewsq ~ L�F&�uq ~ O   q ~�q ~�q ~ gw  �sq ~ '�7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7^xq ~e~q ~e}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ LUZnOuq ~ O   q ~ Qq ~ �q ~7iw  0sq ~ '�9"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~WRxq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~e�sq ~ L;�wuq ~ O   q ~WWw   <sq ~ '�KD�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ L��uq ~ O   q ~&w  0sq ~ 'uւ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
hxq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ L�%SWuq ~ O   q ~
sq ~uw  sq ~ ' &�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~e�sq ~ L ��uq ~ O   q ~�w  
sq ~ 's�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<Lxq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ L�rq�uq ~ O   q ~3q ~ Rw  	#sq ~ '��Gxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t pensacola:nxq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ L^w��uq ~ O   q ~�w  �sq ~ '��|�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8-xq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ LvK��uq ~ O   q ~�q ~�q ~ �w  )sq ~ '��{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ L����uq ~ O   q ~"q ~�w  �sq ~ '�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4xq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~e�sq ~ L��euq ~ O   q ~?q ~+w  �sq ~ '��hAsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~e�q ~e�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fsq ~ L�V3+uq ~ O   q ~Uq ~�w  �sq ~ ''e0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t quincy:nxq ~f
q ~f	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fsq ~ L�u��uq ~ O   q ~�w  �sq ~ '/ҹ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~fq ~fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fsq ~ Lvd�uq ~ O   q ~&�q ~}w  `sq ~ 'KB��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~f&q ~f%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f,sq ~ Lj��uq ~ O   q ~�q ~(�w   sq ~ 'z���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~f3q ~f2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f9sq ~ L�X��uq ~ O   q ~Fq ~ �w  ssq ~ '@�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^�xq ~f@q ~f?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fFsq ~ L╎ uq ~ O   q ~ Qq ~^�w  sq ~ '<�ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t san_antoniot san_antonio:nxq ~fMq ~fLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fVsq ~ L;�uq ~ O   q ~ �q ~)�w  psq ~ '(I sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~M=xq ~f]q ~f\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fcsq ~ Lїuq ~ O   q ~MHq ~xw  Bsq ~ '�X�usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~->xq ~fjq ~fisq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fpsq ~ L�v��uq ~ O   q ~�q ~ w  �sq ~ 'Ѐe�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~fwq ~fvsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f}sq ~ LO�.�uq ~ O   q ~ q ~$q ~"w   �sq ~ 'uk�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_rainiert mount_rainier:mxq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L�Z��uq ~ O   q ~ zt rainierw  �sq ~ '+�ޓsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+rxq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L8��uq ~ O   q ~+}w  sq ~ '��D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L�;�uq ~ O   q ~"q ~"w  �sq ~ 'L���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[�xq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L+(1�uq ~ O   q ~qq ~ w  hsq ~ '.5�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 
mcallen_txt mcallen_tx:cxq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L@��uq ~ O   q ~ Qq ~ �q ~E)w  Wsq ~ '���ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~M_xq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L 5[ruq ~ O   q ~�w  sq ~ '[٫�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L�c�uq ~ O   q ~�q ~�q ~"�w  �sq ~ 'm�S*sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~R�xq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L�Puq ~ O   q ~&zq ~�w  �sq ~ '��	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t clark_fork_rivert clark_fork_river:rxq ~f�q ~f�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~f�sq ~ L?*�uq ~ O   t clarkt forkq ~ �w  @sq ~ '��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~gq ~gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gsq ~ L�8uq ~ O   q ~q ~
q ~�w  �sq ~ '�z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~gq ~gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gsq ~ L*)zVuq ~ O   q ~�q ~ �w  \sq ~ '�_��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bnxq ~gq ~gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g%sq ~ L9��uq ~ O   q ~�q ~*w  
sq ~ '��a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/yxq ~g,q ~g+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g2sq ~ Ly�Fuq ~ O   q ~/�w  Ksq ~ '��V#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~g9q ~g8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g?sq ~ LP��uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  �sq ~ '�{$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0	xq ~gFq ~gEsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gLsq ~ L+�Y�uq ~ O   q ~ Qq ~ �q ~0w  �sq ~ ']��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~gSq ~gRsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gYsq ~ L���uq ~ O   q ~ Qq ~ �q ~hw  �sq ~ ':�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~g`q ~g_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gfsq ~ L�+��uq ~ O   q ~ Qq ~ �q ~ �q ~		w  �sq ~ 's�B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~gmq ~glsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~gssq ~ LR��<uq ~ O   q ~ Rq ~ Sq ~�w   �sq ~ 'pWO�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~gzq ~gysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ LL�O>uq ~ O   q ~Xq ~
�q ~�w  .sq ~ '^���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8|xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L :�uq ~ O   q ~8�w  �sq ~ '�s9[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L��uq ~ O   q ~�q ~ �w  �sq ~ '�L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L{u�uq ~ O   q ~�q ~�w  �sq ~ '�{-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L(k�uq ~ O   q ~ �q ~		q ~ �w  nsq ~ 'E5�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L�C�uq ~ O   q ~ Qq ~�q ~ �w  	�sq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L����uq ~ O   q ~+Vw  	}sq ~ '	��Dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L��vuq ~ O   q ~ Qq ~ �q ~�w  ksq ~ '�p`/sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ LO�Z�uq ~ O   q ~�w  sq ~ 'M6�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t framingham:nxq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~g�sq ~ L���uq ~ O   q ~�w  �sq ~ '5��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~g�q ~g�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hsq ~ Lk\�uq ~ O   q ~ Qq ~ �q ~1w  �sq ~ '3��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~IUxq ~hq ~h
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hsq ~ LTJ=�uq ~ O   q ~�q ~
�q ~�w   sq ~ 'M�.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/4xq ~hq ~hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hsq ~ L��Oquq ~ O   q ~
�q ~�q ~ Rw  �sq ~ 'r���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~G#xq ~h%q ~h$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h+sq ~ L�c�uq ~ O   q ~ Qq ~ �q ~G.w  �sq ~ '_���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~h2q ~h1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h8sq ~ L���Yuq ~ O   q ~,q ~"w  Jsq ~ '�a;qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt west_hartford_ctt west_hartford_ct:cxq ~h?q ~h>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hHsq ~ L�d�uq ~ O   q ~ Qq ~ �q ~q ~Cw  esq ~ ':��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~hOq ~hNsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hUsq ~ Lm�-�uq ~ O   q ~�q ~&cw   sq ~ 'Cg��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~h\q ~h[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hbsq ~ Lw���uq ~ O   q ~ Qq ~ �q ~�w   �sq ~ '[pFWsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ �\� Bt 
<lo,<i,t>>q ~ :q ~Dq ~t population:<lo,<i,t>>xq ~hiq ~hhsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~hssq ~ Ld�wuq ~ O   q ~E"w   =sq ~ '��msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~hzq ~hysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ Lʾ��uq ~ O   q ~
�q ~(�w   �sq ~ 'w��q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~h�q ~h�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~h�sq ~ L ��uq ~ O   t runw  	�sq ~ 'ʨЕsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ L\�#uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t pontchartraint pontchartrain:lxq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ L�SF>uq ~ O   q ~q ~h�w  �sq ~ 'D.�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t west_valleyt west_valley:nxq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ Lբpuq ~ O   q ~q ~w  !sq ~ '���csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4�xq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ LG_��uq ~ O   q ~$q ~$w  �sq ~ '^Om�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Sxq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ L:�+8uq ~ O   q ~ Qq ~ �q ~^w  sq ~ '8)٠q ~Asq ~ sq ~ sq ~ 
w   q ~Eq ~�xq ~h�q ~h�sq ~ @q ~Osq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~h�q ~Xw   ?sq ~ '��Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ L��5puq ~ O   q ~-�q ~ �w  	sq ~ '��U�q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ nt mount_whitneyt mount_whitney:mxq ~h�q ~h�sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~h�sq ~ L+ېuq ~ O   q ~	�w  
+sq ~ '>�*[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t san_bernardinot san_bernardino:nxq ~h�q ~h�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~isq ~ L���6uq ~ O   q ~ �q ~ �w  1sq ~ '4g�qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt richardson_txt richardson_tx:cxq ~iq ~i
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~isq ~ L����uq ~ O   q ~ Qq ~ �q ~O~w  �sq ~ '%�
{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~iq ~isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i!sq ~ L�{��uq ~ O   q ~'q ~5w  	�sq ~ 'X[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~i(q ~i'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i.sq ~ L�qkSuq ~ O   q ~�q ~Aw  Zsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	Exq ~i5q ~i4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i;sq ~ L9��Kuq ~ O   q ~	Pq ~ �q ~�w  sq ~ '�s�q ~sq ~ sq ~ sq ~ 
w   q ~�xq ~iAq ~i@sq ~ @q ~sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~iEq ~w   9sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~iJq ~iIsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~iPsq ~ L�Y�-uq ~ O   q ~<q ~ �w  bsq ~ '�H�asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~iWq ~iVsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i]sq ~ LV��Huq ~ O   q ~�q ~�w  :sq ~ '�j;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
buena_parkt buena_park:nxq ~idq ~icsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~imsq ~ L���uq ~ O   q ~3�q ~pw  	lsq ~ '��g�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~J}xq ~itq ~issq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~izsq ~ L����uq ~ O   q ~gq ~�w  xsq ~ 'NP��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bxq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ LED��uq ~ O   q ~ Qq ~fq ~ �w  �sq ~ '�;��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ Lޟ�{uq ~ O   q ~�q ~�w  <sq ~ 'u0�Sq ~�sq ~ sq ~ sq ~ J   w   q ~Aq ~Hxq ~i�q ~i�sq ~ @q ~�sq ~ G�W9J    sq ~ sq ~ J   w   q ~ �q ~xq ~i�q ~+$w  	�sq ~ '��	psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ Ltcxuq ~ O   q ~�q ~ �w  	Esq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_east_buttresst mount_east_buttress:mxq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ Lɖ`uq ~ O   q ~ zq ~gq ~\�w   sq ~ '6��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t 	atlanta:nxq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ L�NI�uq ~ O   q ~w  	Msq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ L�yIuq ~ O   q ~�w  	3sq ~ 'U1q ~�sq ~ sq ~ sq ~ J   w   q ~xq ~i�q ~i�sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~i�sq ~ L�urIuq ~ O   t citizensw  
sq ~ 'mp�esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6xq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~i�sq ~ L����uq ~ O   q ~
/w  �sq ~ ' 6ƙq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~i�sq ~ L 6NZuq ~ O   t themw  	�sq ~ '5��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~i�q ~i�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jsq ~ L���uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~j
q ~j	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~�xq ~jsq ~ L  �uq ~ O   t now   sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~jq ~jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jsq ~ L�)��uq ~ O   q ~�q ~�w  /sq ~ '˘�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~j%q ~j$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j+sq ~ Lfuq ~ O   q ~ Qq ~ �q ~4w  �sq ~ 'q�S�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Knxq ~j2q ~j1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j8sq ~ L���uq ~ O   q ~,�q ~"w  	sq ~ 'N���q ~�sq ~ sq ~ sq ~ J   w   q ~Mq ~�xq ~j>q ~j=sq ~ @q ~�sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~jBsq ~ L ���uq ~ O   q ~<w  
Csq ~ '�O5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~jIq ~jHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jOsq ~ L9J�Muq ~ O   q ~�q ~"w  -sq ~ '��TXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~?t albany:nxq ~jVq ~jUsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j^sq ~ L��3uq ~ O   q ~?w  }sq ~ '���Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~jeq ~jdsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jksq ~ L��uq ~ O   q ~ Rq ~ Sq ~gw  �sq ~ '�a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t tulsa:nxq ~jrq ~jqsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~jzsq ~ L�y�uq ~ O   q ~�w  �sq ~ '�b�q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~j�q ~jsq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L ���uq ~ O   q ~<w  
Xsq ~ 'e�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t corpus_christit corpus_christi:nxq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ Le��duq ~ O   q ~
q ~
w  sq ~ ']���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L�;�uq ~ O   q ~Uq ~�q ~ Rw  �sq ~ '�G>8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9�xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L���~uq ~ O   q ~
�q ~9�w  �sq ~ ']mCsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L�p*�uq ~ O   q ~6w  �sq ~ 'I�߫sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\Pxq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L�A��uq ~ O   q ~=Oq ~ gw  #sq ~ '鋋sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ LYN�
uq ~ O   q ~ Qq ~ �q ~Nq ~q ~w  tsq ~ '+rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ Lp��7uq ~ O   q ~
�q ~5q ~ �w  �sq ~ '�]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0�xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L���uq ~ O   q ~0�q ~5w  	�sq ~ '�e0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~j�q ~j�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~j�sq ~ L��7�uq ~ O   q ~	�w  dsq ~ 'R���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7@xq ~kq ~ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k	sq ~ L�.}uq ~ O   q ~7Kw  �sq ~ '�Rxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~qt tucson:nxq ~kq ~ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ksq ~ L̑��uq ~ O   q ~qw  ~sq ~ '��!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5�xq ~kq ~ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k%sq ~ L#��uq ~ O   q ~ Qq ~ Rq ~ Sq ~Iw  �sq ~ 'AJ@�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,�xq ~k,q ~k+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k2sq ~ La��"uq ~ O   q ~(�w  �sq ~ '�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~k9q ~k8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k?sq ~ L�Rϻuq ~ O   q ~�q ~_w  	�sq ~ 'G��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bxq ~kFq ~kEsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~kLsq ~ L>��.uq ~ O   q ~fq ~ �w  �sq ~ '�m��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~kSq ~kRsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~kYsq ~ L��uq ~ O   q ~�q ~ Rw  ?sq ~ '�p�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<�xq ~k`q ~k_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~kfsq ~ L�%uq ~ O   q ~�q ~	�w  <sq ~ 'BR�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~kmq ~klsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~kssq ~ L�4�3uq ~ O   q ~'�q ~uw  �sq ~ 'T⭒sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~04xq ~kzq ~kysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L	�9�uq ~ O   q ~0?w  �sq ~ '�ﰹsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	san_diegot san_diego:nxq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L�5huq ~ O   q ~ �q ~�w  xsq ~ '���6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&Xxq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ LG��;uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '� e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L��$�uq ~ O   q ~ q ~	bq ~ w  Fsq ~ '{n:"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L��uq ~ O   q ~Uq ~�w  �sq ~ '�>1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~txq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ LG��uq ~ O   q ~xq ~ Rw  �sq ~ 'J��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_mckinleyt mount_mckinley:mxq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L,�!Muq ~ O   q ~ zt mckinleyw  �sq ~ '_8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7@xq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L��uq ~ O   q ~ Qq ~ �q ~7Kw  sq ~ '�j�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Mt 	spokane:nxq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L�ٲ}uq ~ O   q ~Mw  \sq ~ 'Ԅ0�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$xq ~k�q ~k�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~k�sq ~ L�>D`uq ~ O   q ~�q ~ �w  	sq ~ 'vM{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~lq ~lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lsq ~ LI��5uq ~ O   q ~ Qq ~ �q ~�w  9sq ~ 'ׇ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t tyler:nxq ~lq ~lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lsq ~ L�I�uq ~ O   q ~�w  �sq ~ 'e��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~bjxq ~l!q ~l sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l'sq ~ L��"uq ~ O   q ~ Qq ~buq ~ �w  _sq ~ '�r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t becharoft 
becharof:lxq ~l.q ~l-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l7sq ~ LW�U�uq ~ O   q ~q ~l0w  �sq ~ '%�Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~+}t 	medford:nxq ~l>q ~l=sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lFsq ~ L8��uq ~ O   q ~+}w  usq ~ '�
wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	ann_arbort ann_arbor:nxq ~lMq ~lLsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lVsq ~ L��uq ~ O   q ~*[q ~*\w  �sq ~ '�&�1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~l]q ~l\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lcsq ~ L�f{�uq ~ O   q ~gq ~ Rw  �sq ~ 'U|6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_huntert mount_hunter:mxq ~ljq ~lisq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~lssq ~ Lxo�guq ~ O   q ~ zt hunterw  sq ~ 'l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t davenport:nxq ~l{q ~lzsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ L[���uq ~ O   q ~�w  	csq ~ '��fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t providence:nxq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ L:KMuq ~ O   q ~�w  	:sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
5xq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ Lo3uq ~ O   q ~
@w  �sq ~ '�#�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t bristol_townshipt bristol_township:nxq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ Lߢ�uq ~ O   q ~q ~
w  )sq ~ 'S��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ L!�uq ~ O   q ~Ft wyw  �sq ~ ''^��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ L�<T�uq ~ O   q ~�q ~�w  Csq ~ 'T��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t niagara_fallst niagara_falls:nxq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ LZ
�uq ~ O   q ~�q ~Ew  =sq ~ '�_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~.t 	georgia:nxq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ L�L�uq ~ O   q ~.w  /sq ~ '��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~l�sq ~ L��|~uq ~ O   q ~ q ~w  �sq ~ '�Ҽxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t elizabeth:nxq ~l�q ~l�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~msq ~ L�!@�uq ~ O   q ~�w  .sq ~ '9{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~mq ~msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~msq ~ L�s�uq ~ O   q ~�q ~_w  �sq ~ '��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t irondequoit:nxq ~mq ~msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m!sq ~ L#���uq ~ O   q ~�w  �sq ~ 'e53�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~m(q ~m'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m.sq ~ LX��uq ~ O   q ~ Qq ~�q ~ �w  sq ~ '��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~m5q ~m4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m;sq ~ L�?%uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '5asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ixq ~mBq ~mAsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~mHsq ~ L�dG�uq ~ O   q ~O~q ~w  sq ~ '%Y#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%oxq ~mOq ~mNsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~mUsq ~ L�BA�uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~m\q ~m[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~mbsq ~ Lm�s�uq ~ O   q ~.�w   �sq ~ '�B��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~miq ~mhsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~mosq ~ L�Ȃuq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  /sq ~ '� {psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~mvq ~musq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m|sq ~ L����uq ~ O   q ~&q ~ �w  �sq ~ ',�?�q ~�sq ~ sq ~ sq ~ 
w   q ~Aq ~	!xq ~m�q ~m�sq ~ @q ~�sq ~ G�ǂ    sq ~ sq ~ J   w   q ~ �q ~	,xq ~m�q ~�w   asq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ Lʧ�uq ~ O   q ~ Qq ~ �q ~B�w  Usq ~ 's6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ L}uq ~ O   q ~ Qq ~ Rq ~ Sq ~5w  &sq ~ 'V',�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ L!z�uq ~ O   q ~*q ~ �w  Usq ~ 'W�ڲsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t west_palm_beacht west_palm_beach:nxq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ L����uq ~ O   q ~q ~=q ~	bw  sq ~ '�'D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ LX�7Buq ~ O   q ~3q ~	bw  	1sq ~ '�G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<�xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ L��P;uq ~ O   q ~ Qq ~ �q ~�w  2sq ~ 'j��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ L��Xuq ~ O   q ~ Qq ~ �q ~Hw   �sq ~ '5-�?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ L{\�Vuq ~ O   q ~	�q ~.w  	;sq ~ 'Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~m�q ~m�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~m�sq ~ La�2
uq ~ O   q ~�q ~�q ~�w  �sq ~ '�l{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~nq ~nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n	sq ~ L�V=�uq ~ O   q ~�q ~�w  sq ~ 'cٔ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5xq ~nq ~nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~nsq ~ L��]uq ~ O   q ~S�w   2sq ~ '��gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~nq ~nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n#sq ~ L_uq ~ O   q ~�q ~�w  �sq ~ '<wVsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ Cxq ~n*q ~n)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n0sq ~ L���uq ~ O   q ~ Qq ~ �q ~ Nw  'sq ~ 'R�#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~P�xq ~n7q ~n6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n=sq ~ L[	O�uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w   �sq ~ ' 6Szsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~nDq ~nCsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~nJsq ~ L 5�;uq ~ O   t showw   sq ~ '
�Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_sanfordt mount_sanford:mxq ~nRq ~nQsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n[sq ~ L/�#�uq ~ O   q ~ zt sanfordw  sq ~ '�+�*q ~�sq ~ sq ~ sq ~ J   w   q ~WRxq ~nbq ~nasq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~nfsq ~ L .��uq ~ O   q ~ �w  
Gsq ~ '�TЧsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_massivet mount_massive:mxq ~nmq ~nlsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~nvsq ~ L�kKuq ~ O   q ~ zt massivew  �sq ~ '(�d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0xq ~n~q ~n}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ L�I~2uq ~ O   q ~;w  �sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>�xq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ L�:�uq ~ O   q ~�q ~�q ~�w  �sq ~ '�1Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ L���uq ~ O   q ~ Qq ~ �q ~qw   sq ~ 'R�,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Sxq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ L.���uq ~ O   q ~^w  qsq ~ '�I�Osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~TNxq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ Lt�Suq ~ O   q ~.q ~ Rw   �sq ~ '�"��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~M_xq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ Lv�uq ~ O   q ~�q ~V>w  �sq ~ '�A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~n�sq ~ L���@uq ~ O   q ~!�w   dsq ~ '�&�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~n�sq ~ L��muq ~ O   t whatsw  
'sq ~ '�ߒ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ L��+:uq ~ O   q ~q ~ �w  �sq ~ '�;d;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~n�sq ~ L �~uq ~ O   q ~#q ~(�w  	sq ~ 'S92sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~n�q ~n�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~osq ~ L��t�uq ~ O   q ~=�q ~=�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t new_rochellet new_rochelle:nxq ~o	q ~osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~osq ~ L�&uq ~ O   q ~�q ~#�w  @sq ~ '}w�/q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~oq ~osq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~osq ~ L�k5uq ~ O   t existw  
sq ~ '��q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~o#q ~o"sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~o'sq ~ L  �uq ~ O   t tow  	�sq ~ '�z�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~o/q ~o.sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o5sq ~ Lݯ��uq ~ O   q ~�q ~"w  zsq ~ '"isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Mxq ~o<q ~o;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~oBsq ~ L ���uq ~ O   q ~<w   Xsq ~ 'm�h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@+xq ~oIq ~oHsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~oOsq ~ Lī6duq ~ O   q ~�q ~	�w  Asq ~ 'n��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~{xq ~oVq ~oUsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o\sq ~ L^w��uq ~ O   q ~�w  sq ~ 'Kh��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t el_pasot 	el_paso:nxq ~ocq ~obsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~olsq ~ L 5�&uq ~ O   q ~ �q ~1�w  
sq ~ '+�P[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~osq ~orsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~oysq ~ LQuq ~ O   q ~2�q ~�w  �sq ~ '�#�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~o�sq ~ L�~�Cuq ~ O   t combinedw  
sq ~ 'zպ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~c#xq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ Lj�uq ~ O   q ~ Qq ~c.w  �sq ~ '�q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%�xq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ L?j2�uq ~ O   q ~%5w  psq ~ '�k�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~]zxq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ LOB6Fuq ~ O   q ~ Qq ~ �q ~w   �sq ~ '_��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t tombigbee_rivert tombigbee_river:rxq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ Lm,�uq ~ O   q ~ Qt 	tombigbeew  �sq ~ 'Q�x=sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)xq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ L�9�Guq ~ O   q ~ Qq ~ �q ~)q ~)w  �sq ~ 'x�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ LZ��uq ~ O   q ~2�q ~�w  �sq ~ '"g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_st_eliast mount_st_elias:mxq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ LO��juq ~ O   q ~ zq ~Nt eliasw   �sq ~ '��v�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>xq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ L��)5uq ~ O   q ~>q ~�q ~Fw  �sq ~ 'zH�^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~o�q ~o�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~o�sq ~ Lܠ+.uq ~ O   q ~=�q ~=�q ~"w  }sq ~ 'Q��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ ft 
dearborn:nxq ~pq ~psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~psq ~ LŮ�uq ~ O   q ~ fw  �sq ~ 'e�:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~I}t 	pontiac:nxq ~pq ~psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~psq ~ L�hDduq ~ O   q ~I}w  �sq ~ 'R��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~$�t cleveland:nxq ~p$q ~p#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p,sq ~ L�h�tuq ~ O   q ~$�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;;xq ~p3q ~p2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p9sq ~ L�$u�uq ~ O   q ~;Fq ~q ~"w  jsq ~ '��4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt fort_worth_txt fort_worth_tx:cxq ~p@q ~p?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~pIsq ~ L��uq ~ O   q ~ �q ~CCw  Xsq ~ '�CQsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@�xq ~pPq ~pOsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~pVsq ~ L��uq ~ O   q ~@�w  �sq ~ '�}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~p]q ~p\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~pcsq ~ L�B;uq ~ O   q ~ Qq ~ �q ~w  csq ~ 'U��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Ixq ~pjq ~pisq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ppsq ~ L�B�Duq ~ O   q ~1�w  _sq ~ '��Uxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	abilene:nxq ~pwq ~pvsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~psq ~ L�q��uq ~ O   q ~�w  sq ~ '\�o�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ L��o�uq ~ O   q ~ Qq ~ �q ~"	w  �sq ~ '*l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t great_fallst great_falls:nxq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ L�Kuq ~ O   q ~Dq ~Ew  �sq ~ '��b�q ~�sq ~ q ~Swq ~Swsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~p�q ~Q�w  	�sq ~ '�ZQ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&ixq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ L��:uq ~ O   q ~�q ~ �w  �sq ~ 'fI��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ L��5uq ~ O   q ~Gw  ]sq ~ '��I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ L�[Guq ~ O   q ~)q ~xw  ysq ~ '�e3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ L�Y{uq ~ O   q ~�w  sq ~ '��P�q ~	sq ~ sq ~ sq ~ 
w   q ~�xq ~p�q ~p�sq ~ @q ~	'sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~p�q ~	.w    sq ~ '�YS�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~p�sq ~ L�Xۇuq ~ O   t numberw  
-sq ~ 'OG�q ~�sq ~ sq ~ sq ~ 
w   q ~Axq ~p�q ~p�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~p�q ~�w   sq ~ '-R��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<xq ~p�q ~p�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~p�sq ~ Laz�uq ~ O   q ~Gq ~ �w  �sq ~ '⏩�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t simi_valleyt simi_valley:nxq ~qq ~qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qsq ~ L�kouq ~ O   q ~;Fq ~w  �sq ~ 'ċz�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~qq ~qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qsq ~ L�b!kuq ~ O   q ~7q ~w  �sq ~ 'w�\fq ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~qq ~qsq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~q#sq ~ L 0luq ~ O   t floww  
!sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<Lxq ~q+q ~q*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q1sq ~ L8�quq ~ O   q ~3w  xsq ~ '�x��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3�xq ~q8q ~q7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q>sq ~ L���uq ~ O   q ~3�q ~pw  �sq ~ '��ݙsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~qEq ~qDsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qKsq ~ L5<_uq ~ O   q ~Dq ~Eq ~�w  Usq ~ ':���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~qRq ~qQsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qXsq ~ L�C�7uq ~ O   q ~	�q ~�w  �sq ~ '��#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q_q ~q^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qesq ~ LӺuq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
Fxq ~qlq ~qksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qrsq ~ L^[ީuq ~ O   q ~
Qq ~+Vw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~qyq ~qxsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~qsq ~ L���#uq ~ O   q ~q ~=w  $sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0Exq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L����uq ~ O   q ~<q ~=w  �sq ~ '��L�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ LON��uq ~ O   q ~�q ~�q ~�w  |sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)�xq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L�.�uq ~ O   q ~ �q ~)�q ~w  sq ~ '(�?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~;t bloomington:nxq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L�I~2uq ~ O   q ~;w  sq ~ '߰~4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~D�xq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L �{|uq ~ O   q ~D�q ~D�w  �sq ~ '���<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L�J�(uq ~ O   q ~ Qq ~�w  �sq ~ '`�R�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L16�uq ~ O   q ~�w   �sq ~ '���q ~]sq ~ sq ~ sq ~ 
w   q ~Hxq ~q�q ~q�sq ~ @q ~]sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~q�q ~]w   sq ~ 'e��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0Exq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L:�>Fuq ~ O   q ~<q ~ w  �sq ~ '~6� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bnxq ~q�q ~q�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~q�sq ~ L3�IKuq ~ O   q ~�q ~xw  �sq ~ '�Ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~rq ~rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~rsq ~ L�W%uq ~ O   q ~Ww  �sq ~ '#{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~rq ~rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~rsq ~ L�
uq ~ O   q ~Fq ~�w  sq ~ '��%;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'axq ~rq ~rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r%sq ~ L��6uq ~ O   q ~'lq ~w  �sq ~ '��}xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ �t elyria:nxq ~r,q ~r+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r4sq ~ L��Vuq ~ O   q ~ �w  /sq ~ 'υ9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~r;q ~r:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~rAsq ~ L-tpwuq ~ O   q ~Dq ~w  sq ~ '&�:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t santa_monicat santa_monica:nxq ~rHq ~rGsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~rQsq ~ L��.uq ~ O   q ~ q ~;w  �sq ~ '!��=sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~f�xq ~rXq ~rWsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r^sq ~ L4��ruq ~ O   q ~E)w  �sq ~ '��n8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ ��zPt <s,c>q ~ 8q ~ Zq ~<t capital:<s,c>xq ~req ~rdsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~rosq ~ L ���uq ~ O   q ~<w   8sq ~ '�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~G.t 
mesquite:nxq ~rvq ~rusq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r~sq ~ L�a�9uq ~ O   q ~G.w  tsq ~ 'r� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L�ץuuq ~ O   q ~ Qq ~ �q ~Gw  Fsq ~ 'Ujsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;�xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L�P�uq ~ O   q ~3sq ~Uw  �sq ~ '¸�4sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'rxq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L8�auq ~ O   q ~'}q ~w  Msq ~ 'ߚ�Asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L����uq ~ O   q ~ Rq ~ Sq ~�q ~�w  �sq ~ '�ҝhsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L���uq ~ O   q ~Wq ~!�w  sq ~ '+{�Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L�D�Luq ~ O   q ~ Qq ~ �q ~�w  Lsq ~ 'lN=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3�xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ L(�Auq ~ O   q ~ Qq ~ �q ~3�q ~pw  sq ~ 'k1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,{xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ Lq0ouq ~ O   q ~'0q ~"w  �sq ~ '��Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~r�sq ~ LrB�uq ~ O   q ~ Qq ~ Rq ~ Sq ~Uq ~
�w  �sq ~ '�׀sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~r�q ~r�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s sq ~ L���uq ~ O   q ~Dw  �sq ~ '��rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~sq ~ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ssq ~ L0fBuq ~ O   q ~ Qq ~ �q ~=�q ~=�w  �sq ~ '��Y�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t champaign:nxq ~sq ~ssq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ssq ~ LU��uq ~ O   q ~�w  �sq ~ 'ۧg{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~s#q ~s"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s)sq ~ L�ץ1uq ~ O   q ~
�w  �sq ~ '��Ԕq ~�sq ~ sq ~ sq ~ J   w   q ~xq ~s/q ~s.sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~s3q ~	w  	�sq ~ 'a��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Ixq ~s8q ~s7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s>sq ~ L�{;�uq ~ O   q ~ Qq ~ �q ~1�w  >sq ~ 't��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t st_clair_shorest st_clair_shores:nxq ~sEq ~sDsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sNsq ~ Lyp�$uq ~ O   q ~Nq ~q ~w  wsq ~ 'ab��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/	xq ~sUq ~sTsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s[sq ~ L?�#�uq ~ O   q ~ Qq ~ �q ~/w  Bsq ~ 'r�)ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~sbq ~sasq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~shsq ~ L��W�uq ~ O   q ~ Qq ~ �q ~L�q ~ �w  �sq ~ ' `\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~soq ~snsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~susq ~ L�uq ~ O   q ~ Qq ~8�w  	Tsq ~ 'w���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~s|q ~s{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~s�sq ~ L ��uq ~ O   q ~w   Jsq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~s�sq ~ L z�uq ~ O   q ~`'w   sq ~ '�?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"sxq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L/�+uq ~ O   q ~�w  	fsq ~ 'SN�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L|�`�uq ~ O   q ~#q ~ �w  �sq ~ '��{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'}t erie:nxq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L /��uq ~ O   q ~'}w   sq ~ '�R�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~?axq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L��7uq ~ O   q ~8�q ~0�w  Ssq ~ 'K��Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
Fxq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L���huq ~ O   q ~
Qw  �sq ~ 'J��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L��:uq ~ O   q ~gq ~hq ~�q ~Fw  �sq ~ ',O��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_quandaryt mount_quandary:mxq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ Ls�K<uq ~ O   q ~ zt quandaryw  Psq ~ '�u��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~s�q ~s�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~s�sq ~ L�X��uq ~ O   q ~ Qq ~ �q ~�q ~	bw  �sq ~ '!�f�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
maryland:nxq ~tq ~tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tsq ~ L���uq ~ O   q ~�w  �sq ~ '[���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~tq ~tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tsq ~ L8$�uq ~ O   q ~Xq ~�w  Vsq ~ '�H�:sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~F#xq ~t q ~tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t&sq ~ L���*uq ~ O   q ~ Qq ~ �q ~F.w  ~sq ~ '�*�q ~=sq ~ sq ~ sq ~ 
w   q ~Aq ~Hxq ~t,q ~t+sq ~ @q ~Lsq ~ G�W9J    sq ~ sq ~ J   w   q ~ �q ~xq ~t0q ~Qw   fsq ~ '���)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8Mxq ~t5q ~t4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t;sq ~ Lk�RDuq ~ O   q ~8Xq ~ �w  sq ~ ' v�Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2xq ~tBq ~tAsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tHsq ~ L�s�1uq ~ O   q ~ zq ~�w  sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Dt allentown:nxq ~tOq ~tNsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tWsq ~ L���uq ~ O   q ~Dw  �sq ~ 'n��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"�xq ~t^q ~t]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tdsq ~ L����uq ~ O   q ~
/w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~tkq ~tjsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~tqsq ~ L��uq ~ O   q ~
�q ~w   �sq ~ '�L�#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~txq ~txq ~twsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t~sq ~ LT�� uq ~ O   q ~ Qq ~ Rq ~ Sq ~xw  ]sq ~ '�i�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_princetont mount_princeton:mxq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ LTO�Quq ~ O   q ~ zt 	princetonw  �sq ~ 'm�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ LP�-uq ~ O   q ~Nq ~q ~q ~ gw  %sq ~ '�)Lq ~-sq ~ sq ~ sq ~ 
w   q ~	!xq ~t�q ~t�sq ~ @q ~-sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~t�q ~-w   Ssq ~ '��͢sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ L�h��uq ~ O   q ~qq ~B�w  	�sq ~ '��JBsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ L��61uq ~ O   q ~�q ~B�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'?xq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ L���uq ~ O   q ~'Jq ~0�w  �sq ~ 'Y	:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
fort_smitht fort_smith:nxq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ LYDxuq ~ O   q ~ �q ~ �w  Jsq ~ '?�jpsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~pAxq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ L���?uq ~ O   q ~ �q ~CCq ~w  �sq ~ '>��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~<t 	roanoke:nxq ~t�q ~t�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~t�sq ~ LQz��uq ~ O   q ~<w  hsq ~ '\o�<q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~t�sq ~ L\o�uq ~ O   t runningw  	�sq ~ 'U*��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/	xq ~uq ~usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~usq ~ L3O��uq ~ O   q ~/w  usq ~ '�:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~uq ~usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~usq ~ LLɅpuq ~ O   q ~ Qq ~ �q ~�w   �sq ~ '��y?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~u!q ~u sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u'sq ~ L:ɂuq ~ O   q ~ Qq ~ �q ~w  @sq ~ '��x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~TNxq ~u.q ~u-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u4sq ~ L�:�uq ~ O   q ~ Rq ~ Sq ~.w  	`sq ~ '�Y�Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~_xq ~u;q ~u:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~uAsq ~ LΫuq ~ O   q ~ Qq ~ Rq ~ Sq ~iw  -sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~uHq ~uGsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~uNsq ~ L�w��uq ~ O   q ~�q ~(�w  �sq ~ 'y݋!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t grand_prairiet grand_prairie:nxq ~uUq ~uTsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u^sq ~ L�#xuq ~ O   q ~�q ~�w  �sq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$xq ~ueq ~udsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~uksq ~ L�20Buq ~ O   q ~ Qq ~ �q ~�w  Esq ~ '"2��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~:xq ~urq ~uqsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~uxsq ~ L�k^�uq ~ O   q ~Eq ~(�w  	0sq ~ 'dà�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_vancouvert mount_vancouver:mxq ~uq ~u~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ L�`�Duq ~ O   q ~ zt 	vancouverw  &sq ~ 'm|��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~vxq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ LR��]uq ~ O   q ~ Qq ~ �q ~�w  	�sq ~ '6I'Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ L-uuq ~ O   q ~*q ~"w  	sq ~ 'B��?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Eq ~	!xq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~u�sq ~ L 3;�uq ~ O   q ~w   csq ~ ',�"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
hxq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ L�{��uq ~ O   q ~ Qq ~ �q ~
sw  �sq ~ '��V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ L��,tuq ~ O   q ~�q ~�w   �sq ~ '�8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	!xq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~u�sq ~ LW��uq ~ O   q ~ Qq ~	0w   Bsq ~ 'ȴKLsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Dxq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ L��t�uq ~ O   q ~�q ~3w  Gsq ~ 'G�X�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~!�t 	reading:nxq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~u�sq ~ L@e��uq ~ O   q ~!�w  Dsq ~ '8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t flatheadt 
flathead:lxq ~u�q ~u�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vsq ~ Lg
uq ~ O   q ~q ~u�w  �sq ~ '-I|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>�xq ~v
q ~v	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vsq ~ Lz	�uq ~ O   q ~ Qq ~>�w   �sq ~ 'W@�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~vq ~vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vsq ~ L]�w�uq ~ O   q ~gq ~/q ~0q ~ �w  �sq ~ 'D��Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t dearborn_heightst dearborn_heights:nxq ~v$q ~v#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v-sq ~ L����uq ~ O   q ~ fq ~�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t iliamnat 	iliamna:lxq ~v4q ~v3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v=sq ~ Lvη�uq ~ O   q ~q ~v6w  ksq ~ 'h���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~->xq ~vDq ~vCsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vJsq ~ Lv�y:uq ~ O   q ~�q ~=w  �sq ~ '��e{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t oak_lawnt 
oak_lawn:nxq ~vQq ~vPsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vZsq ~ L f�3uq ~ O   q ~�q ~	sw  �sq ~ '{Zܥsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+rxq ~vaq ~v`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vgsq ~ L����uq ~ O   q ~+}q ~�w  �sq ~ '�"��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~vnq ~vmsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~vtsq ~ L�<�uq ~ O   q ~ Qq ~ �q ~�w  	�sq ~ '�n xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	concord:nxq ~v{q ~vzsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ L8��^uq ~ O   q ~�w  �sq ~ 'L~Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t superiort 
superior:lxq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ L�cV�uq ~ O   q ~q ~v�w  �sq ~ 'x�J�q ~nsq ~ sq ~ sq ~ 
w   q ~�q ~5xq ~v�q ~v�sq ~ @q ~nsq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~v�q ~nw   Osq ~ '
ĳ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ L��8uq ~ O   q ~+Ft kyw  �sq ~ '%W��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ gt 
michigan:nxq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ L�)�uq ~ O   q ~ gw  ,sq ~ '\�+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
okeechobeet okeechobee:lxq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ LtnEuq ~ O   q ~q ~v�w  �sq ~ 'z{esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ L�Ы�uq ~ O   q ~Gq ~�w  �sq ~ '��Y;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Knxq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ L��uq ~ O   q ~,�q ~ �w  6sq ~ '��kq ~�sq ~ sq ~ sq ~ J   w   q ~5cxq ~v�q ~v�sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ LY�!+uq ~ O   q ~�w  	�sq ~ '�5\qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~v�q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~v�sq ~ LΏ{uq ~ O   q ~q ~ Rw  sq ~ 'v�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t iowa:nxq ~w q ~v�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wsq ~ L 1j�uq ~ O   q ~�w   �sq ~ 'D��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~wq ~wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wsq ~ L���uq ~ O   q ~. w   �sq ~ '�
�ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	new_havent new_haven:nxq ~wq ~wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w%sq ~ L�Fuq ~ O   q ~�q ~�w  Asq ~ '�)�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t oregon:nxq ~w,q ~w+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w4sq ~ L��ޢuq ~ O   q ~�w  Qsq ~ 't�J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~f�xq ~w;q ~w:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wAsq ~ L�*uq ~ O   q ~ Qq ~f�q ~g q ~ �w  �sq ~ 'Bw�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~txq ~wHq ~wGsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wNsq ~ L��Suuq ~ O   q ~xw  �sq ~ '��R?sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~wUq ~wTsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w[sq ~ L C��uq ~ O   q ~I�q ~.w  	tsq ~ '\(c�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~dxq ~wbq ~wasq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~whsq ~ Lp��uq ~ O   q ~ Qq ~Nq ~d&q ~ �w  2sq ~ '�6]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7�xq ~woq ~wnsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~wusq ~ Lh!��uq ~ O   q ~ Qq ~ �q ~7�w  �sq ~ '0H6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~w|q ~w{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L���uq ~ O   q ~�w  �sq ~ '?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~?�xq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L"��muq ~ O   q ~?�w  �sq ~ 'R�Q)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Knxq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ Lۈ��uq ~ O   q ~ Qq ~ �q ~,�w  .sq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~	�t newark:nxq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L�{��uq ~ O   q ~	�w   �sq ~ '��x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%Qxq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L���Quq ~ O   q ~%\q ~�w  	�sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L�S3uuq ~ O   q ~ Qq ~ �q ~&w  	sq ~ '{`�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%	xq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L��uq ~ O   q ~%w  ,sq ~ 'p�L8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t scottsdale:nxq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L�߲huq ~ O   q ~�w  hsq ~ '�N��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>xq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L�Lq�uq ~ O   q ~>w  (sq ~ '�!*sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~P�xq ~w�q ~w�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~w�sq ~ L�גuq ~ O   q ~�q ~ Rw  !sq ~ ' 0g1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'axq ~xq ~xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xsq ~ L[9,uq ~ O   q ~'lw  Vsq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
Qt anchorage:nxq ~xq ~xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xsq ~ L���huq ~ O   q ~
Qw  sq ~ '��Fq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~xsq ~ L���@uq ~ O   q ~!�w  
_sq ~ '|�'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\�xq ~x&q ~x%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x,sq ~ LW�uq ~ O   q ~\�q ~�w  {sq ~ 'E�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~drxq ~x3q ~x2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x9sq ~ L��B�uq ~ O   q ~�w  �sq ~ 'Rma�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
missouri:nxq ~x@q ~x?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xHsq ~ L���uq ~ O   q ~�w  �sq ~ '\���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t new_bedfordt new_bedford:nxq ~xOq ~xNsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xXsq ~ L�`��uq ~ O   q ~�q ~.w  Psq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ht orange:nxq ~x_q ~x^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xgsq ~ L��&luq ~ O   q ~hw  sq ~ 'll��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*Axq ~xnq ~xmsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xtsq ~ Lأ{�uq ~ O   q ~ Rq ~ Sq ~�w  asq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'[t 	hammond:nxq ~x{q ~xzsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ L)Ac�uq ~ O   q ~'[w  �sq ~ '̇0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>xq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ Lۄ�Kuq ~ O   q ~ Qq ~ �q ~>w   sq ~ '��Uysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	san_mateot san_mateo:nxq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ Lc�
uq ~ O   q ~ �q ~$zw  �sq ~ 'N�Ƹsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t knoxville:nxq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ L^��uq ~ O   q ~�w  ,sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
fort_waynet fort_wayne:nxq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ L�i[uq ~ O   q ~ �q ~�w  �sq ~ '��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~x�sq ~ L�a�uq ~ O   q ~Zw  
sq ~ 'ʬњq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~x�sq ~ LʬY[uq ~ O   t squarew  	�sq ~ '�e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t cedar_rapidst cedar_rapids:nxq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ Lv��Duq ~ O   q ~�q ~�w  	8sq ~ '�k�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_shastat mount_shasta:mxq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ L�w��uq ~ O   q ~ zt shastaw  sq ~ '�쉛sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~x�q ~x�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~x�sq ~ Lr4�Iuq ~ O   q ~Uq ~
�w  �sq ~ '0]��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~yq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ysq ~ LcZ�6uq ~ O   q ~q ~ w  Bsq ~ '=W�Bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~exq ~yq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ysq ~ Lj��uq ~ O   q ~ Qq ~ �q ~pw  �sq ~ '�	��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Irxq ~yq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y%sq ~ L�hDduq ~ O   q ~I}w  �sq ~ '�_H#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~afxq ~y,q ~y+sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y2sq ~ L�(�uq ~ O   q ~ Qq ~ Rq ~ Sq ~}w  [sq ~ '��A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ �t texas:nxq ~y9q ~y8sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~yAsq ~ L�^�uq ~ O   q ~ �w  �sq ~ '�}[xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~P�xq ~yHq ~yGsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~yNsq ~ L 4�uq ~ O   q ~�w  Tsq ~ 'c��]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\Pxq ~yUq ~yTsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y[sq ~ L ͎uq ~ O   q ~=Ow  4sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~J}xq ~ybq ~yasq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~yhsq ~ L�~^�uq ~ O   q ~gq ~w  msq ~ '^ƛ6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~yoq ~ynsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~yusq ~ L��b�uq ~ O   q ~Hw  �sq ~ 'S��Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~y|q ~y{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L3��&uq ~ O   q ~+�q ~w  �sq ~ '��@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/�xq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L~��uq ~ O   q ~/�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&xq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L�Dn�uq ~ O   q ~&w  �sq ~ 'H��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L��~�uq ~ O   q ~ Rq ~ Sq ~�w  sq ~ '�1�=sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L\%�zuq ~ O   q ~ Qq ~ �q ~+Fw  sq ~ 'Xu�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_elbertt mount_elbert:mxq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ Lr���uq ~ O   q ~ zt elbertw  lsq ~ '�'R8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
st greenwich:nxq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L{CDxuq ~ O   q ~
sw  Hsq ~ '�eV�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t fresno:nxq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L��m�uq ~ O   q ~�w   �sq ~ '�u�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7yxq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~y�sq ~ L�0y�uq ~ O   q ~7�q ~ gw  	�sq ~ 'ݐ�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_el_dientet mount_el_diente:mxq ~y�q ~y�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~zsq ~ L��mouq ~ O   q ~ zq ~ �t dientew  �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
@t 	salinas:nxq ~z
q ~z	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~zsq ~ Lo3uq ~ O   q ~
@w  sq ~ '6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~%t dallas:nxq ~zq ~zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z!sq ~ L�.?�uq ~ O   q ~%w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~z(q ~z'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z.sq ~ L;Ro�uq ~ O   q ~ Qq ~ �q ~�q ~�w  	Ysq ~ '�c7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~z5q ~z4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z;sq ~ Ls��uq ~ O   q ~ Qq ~ �q ~Tw  	$sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~zBq ~zAsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~zHsq ~ L��uq ~ O   q ~ Qq ~ �q ~
�w  	Xsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~+�t pomona:nxq ~zOq ~zNsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~zWsq ~ L�n1�uq ~ O   q ~+�w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;�xq ~z^q ~z]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~zdsq ~ LB��cuq ~ O   q ~3sq ~5w  �sq ~ '�	UQsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t baton_rouget baton_rouge:nxq ~zkq ~zjsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ztsq ~ L�B�buq ~ O   q ~�q ~�w  ssq ~ '�]Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\�xq ~z{q ~zzsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L�z�9uq ~ O   q ~\�w  ]sq ~ '�c(�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Zt 	irving_txt irving_tx:cxq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L{��uq ~ O   q ~?�q ~w  �sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~z�sq ~ L  huq ~ O   t isw   sq ~ 'j#sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L��u�uq ~ O   q ~
q ~�w  Jsq ~ 'V��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t peoria:nxq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L��9�uq ~ O   q ~�w   �sq ~ 'J���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ LE��uq ~ O   q ~�q ~�q ~ Rw  Osq ~ '9�%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~z�xq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L����uq ~ O   q ~ Qq ~ �q ~?�w  �sq ~ '%3��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L�*2uq ~ O   q ~2�q ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L?���uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  8sq ~ '�E?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~afxq ~z�q ~z�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~z�sq ~ L� �uq ~ O   q ~}q ~ Rw  	Qsq ~ 'T��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~{q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{	sq ~ L�n1�uq ~ O   q ~+�w  �sq ~ 'o`�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!uxq ~{q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{sq ~ L~D�uq ~ O   q ~ Qq ~ �q ~ �q ~!�w  dsq ~ ' /��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~{q ~{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~{#sq ~ L /"�uq ~ O   t doesw   sq ~ '���\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~{+q ~{*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{1sq ~ L�hO�uq ~ O   q ~aw  	&sq ~ '`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~MNxq ~{8q ~{7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{>sq ~ L%��5uq ~ O   q ~MYq ~ �w  Osq ~ '�]V�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~{Fsq ~ L�\�[uq ~ O   t averagew  	�sq ~ '-g֒sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	6xq ~{Nq ~{Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{Tsq ~ L��6�uq ~ O   q ~ Rq ~ Sq ~�w  �sq ~ 'ͥ,�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~{[q ~{Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{asq ~ L{�"�uq ~ O   q ~Fq ~Uw   �sq ~ 'eP|�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1�xq ~{hq ~{gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{nsq ~ L{��uq ~ O   q ~ Qq ~ �q ~ �q ~1�w  sq ~ '�Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[�xq ~{uq ~{tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{{sq ~ LΉ�Wuq ~ O   q ~qq ~=w  �sq ~ ':��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L%�Wuq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�8n�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~18xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L�uq ~ O   q ~1Cw  Hsq ~ '��Jksq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	teshekpukt teshekpuk:lxq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L���uq ~ O   q ~q ~{�w  sq ~ 'D@��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L��Ғuq ~ O   q ~�q ~�w  �sq ~ 'T LIsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ LB���uq ~ O   q ~2�w  �sq ~ 'ћx�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~K�xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L[�Yuq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  �sq ~ 'C���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L�3T�uq ~ O   q ~ �q ~�w  �sq ~ '4>J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~&�t joliet:nxq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L�0��uq ~ O   q ~&�w  msq ~ '��
�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$oxq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~{�sq ~ L�9:duq ~ O   q ~ Qq ~ �q ~ �q ~$zw  ?sq ~ 'I�t�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)�xq ~{�q ~{�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|sq ~ L��Guq ~ O   q ~ q ~/Lw  	sq ~ 'k�l[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ixq ~|	q ~|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|sq ~ L��(�uq ~ O   q ~ Qq ~ �q ~�q ~tw  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
t wilmington:nxq ~|q ~|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|sq ~ Lp��uq ~ O   q ~
w  `sq ~ '�(��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~|%q ~|$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|+sq ~ L9��9uq ~ O   q ~�q ~ w  	)sq ~ 'Ҵɸsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	houston:nxq ~|2q ~|1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|:sq ~ LA�Ōuq ~ O   q ~�w  asq ~ 'cY�isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~|Aq ~|@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|Gsq ~ L��C�uq ~ O   q ~#q ~�q ~Fw  �sq ~ 'Vh�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt 
mount_beart mount_bear:mxq ~|Nq ~|Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|Wsq ~ L��^�uq ~ O   q ~ zt bearw  �sq ~ 'WmAsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0�xq ~|_q ~|^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|esq ~ L=��uq ~ O   q ~ q ~ Rw  	�sq ~ 'S��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~|lq ~|ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|rsq ~ Lq�uq ~ O   q ~Hq ~ gw   qsq ~ '��
q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~|zsq ~ L�#�uq ~ O   t aboutw  	�sq ~ '��jq ~�sq ~ sq ~ sq ~ J   w   q ~xq ~|�q ~|�sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~|�sq ~ L 6�uq ~ O   t stayw  
Psq ~ '�@��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7 xq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ L�d�4uq ~ O   q ~ Qq ~ �q ~�w  ;sq ~ '��q ~�sq ~ sq ~ sq ~ J   w   q ~5xq ~|�q ~|�sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~|�sq ~ L }>uq ~ O   q ~�w  	�sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Dxq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ Lw�suq ~ O   q ~�q ~~w  	-sq ~ 'A���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~pAxq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ L�hI]uq ~ O   q ~ Qq ~ �q ~ �q ~CCw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\zxq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ LC+Muq ~ O   q ~_q ~-�w  csq ~ '�m(;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ L��nuq ~ O   q ~&�q ~w  �sq ~ '�s��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@+xq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ L���uq ~ O   q ~ Qq ~ �q ~�w  Zsq ~ 'f{]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~G#xq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ L�a�9uq ~ O   q ~G.w  �sq ~ 'x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~|�sq ~ L\Uh!uq ~ O   q ~�q ~ �w  �sq ~ 'x�B&sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~|�q ~|�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}sq ~ L�W`uq ~ O   q ~ Qq ~ �q ~w  �sq ~ '�aXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4�xq ~}q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}sq ~ L��uuq ~ O   q ~$q ~$q ~&cw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7^xq ~}q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}sq ~ LI!��uq ~ O   q ~7iw  &sq ~ '* �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Bxq ~}&q ~}%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~},sq ~ L�\�Kuq ~ O   q ~Mq ~�w  �sq ~ 'b�.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~]xq ~}3q ~}2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}9sq ~ L 0L�uq ~ O   q ~hw  ssq ~ 'm�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~}@q ~}?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}Fsq ~ Li�Euq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '4 ;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	st_josepht st_joseph:nxq ~}Mq ~}Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}Vsq ~ L�5t.uq ~ O   q ~Nq ~�w  sq ~ '�zm;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,�xq ~}]q ~}\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}csq ~ L��uq ~ O   q ~(�q ~ �w  esq ~ '�5�6q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~}iq ~}hsq ~ @q ~�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~}mq ~�w   @sq ~ '�ޥ;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'rxq ~}rq ~}qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}xsq ~ L��huq ~ O   q ~'}q ~�w  4sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~}q ~}~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L�	��uq ~ O   q ~ Qq ~ �q ~�w  \sq ~ ')�O�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t arlington_heightst arlington_heights:nxq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L+@uq ~ O   q ~�q ~�w  �sq ~ 'z�9jq ~B�sq ~ sq ~ sq ~ 
w   q ~�xq ~}�q ~}�sq ~ @q ~B�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~}�q ~B�w   sq ~ '���gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L�>uq ~ O   q ~)w   �sq ~ '�Q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<�xq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L�yicuq ~ O   q ~ Qq ~ �q ~<�w  	sq ~ '�K��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"-xq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L�ܾuq ~ O   q ~ Qq ~ �q ~{w  sq ~ '�ߚ1sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L��Yuq ~ O   q ~ Qq ~ �q ~ q ~	bw  sq ~ '2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L�Y5�uq ~ O   q ~#q ~B�q ~Aw   �sq ~ 'g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Gt fairfield:nxq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L�[��uq ~ O   q ~Gw  usq ~ '�B-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Irxq ~}�q ~}�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~}�sq ~ L����uq ~ O   q ~ Qq ~ �q ~I}w  qsq ~ 't�fXq ~�sq ~ sq ~ sq ~ J   w   q ~;xq ~~ q ~}�sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~~sq ~ L ���uq ~ O   q ~<w  	�sq ~ 'X	��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~+�xq ~~q ~~
sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~sq ~ L�z�uq ~ O   q ~+�q ~"w   �sq ~ '�2Ygsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~h�xq ~~q ~~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~sq ~ L��Muq ~ O   q ~ zq ~>xw  Zsq ~ '����q ~�sq ~ q ~Swq ~Swsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~~&q ~x�w  
 sq ~ '�-��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~~+q ~~*sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~1sq ~ L���uq ~ O   q ~hq ~ �w  �sq ~ '�s�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
hxq ~~8q ~~7sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~>sq ~ L{CDxuq ~ O   q ~
sw  ssq ~ '�䑽sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#�xq ~~Eq ~~Dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~Ksq ~ LH�quq ~ O   q ~#�q ~ �w  �sq ~ 'w��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~~Rq ~~Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~~Xsq ~ L 0��uq ~ O   q ~w   *sq ~ '�h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~~_q ~~^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~esq ~ L��uq ~ O   q ~ Rq ~ Sq ~Uq ~�w  Hsq ~ '��8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~~lq ~~ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~rsq ~ LŢ��uq ~ O   q ~�q ~�w  	�sq ~ '��usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~~yq ~~xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~sq ~ L�҉�uq ~ O   q ~�q ~?�w  �sq ~ '�?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t newport_beacht newport_beach:nxq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ LX�7Buq ~ O   q ~3q ~	bw  �sq ~ '�~[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"=xq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ L����uq ~ O   q ~�q ~ �w  qsq ~ 'sʇsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"exq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ LZ�Jbuq ~ O   q ~?q ~�q ~�w  rsq ~ '%�qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~IUxq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ LF��Auq ~ O   q ~�q ~?�w  *sq ~ '��ۑsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	yxq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ L�{��uq ~ O   q ~	�w  �sq ~ '��>q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~~�sq ~ L�P�uq ~ O   t couldw  
9sq ~ '�b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~_xq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ Lm��uq ~ O   q ~iq ~ Rw  
sq ~ '�J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<�xq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ L�@��uq ~ O   q ~<�w   �sq ~ '��d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~~�q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~~�sq ~ L|���uq ~ O   q ~�q ~�q ~_w  >sq ~ '��M�q ~�sq ~ q ~Swq ~Swsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~~�q ~{Gw  	�sq ~ '�7�Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~ q ~~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LƤ��uq ~ O   q ~ Qq ~ Rq ~ Sq ~Sw  csq ~ 'x��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t rochester:nxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L=b�uq ~ O   q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~B�xq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~"sq ~ L���uq ~ O   q ~#q ~B�q ~#w  �sq ~ '3� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Q\xq ~)q ~(sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~/sq ~ L�jO�uq ~ O   q ~ Qq ~ �q ~Fw  esq ~ 'P��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~_t 
portland:nxq ~6q ~5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~>sq ~ L+u*uq ~ O   q ~_w  sq ~ 'A�r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Eq ~Dsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~Ksq ~ Lz�p�uq ~ O   t sparsestw   sq ~ 'k��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~}xq ~Sq ~Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Ysq ~ L 6u&uq ~ O   q ~�w  �sq ~ '��Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~`q ~_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~fsq ~ Lz��6uq ~ O   q ~ Qq ~ Rq ~ Sq ~
�q ~
�w  hsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)wxq ~mq ~lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ssq ~ L�轇uq ~ O   q ~�q ~�q ~ �w  �sq ~ ''\��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Q\xq ~zq ~ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�1�Kuq ~ O   q ~Fw  �sq ~ '�d��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LD��uq ~ O   q ~ Qq ~ �q ~�w  sq ~ 'փ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~P�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�{Vquq ~ O   q ~B�q ~ Rw   xsq ~ ':�Uxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
billings:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L5-�uq ~ O   q ~�w  	Hsq ~ '�ƐCsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�+]uq ~ O   q ~�q ~Uw  �sq ~ 'Bl0�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~&�t waco:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L 7��uq ~ O   q ~&�w  �sq ~ 'ɒV[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lz��uq ~ O   q ~q ~+w  hsq ~ '�<�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~h@xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�?�huq ~ O   q ~q ~Cq ~uw  esq ~ '�?J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Kxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LI�љuq ~ O   q ~Vq ~"�w  �sq ~ '��f�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_lincolnt mount_lincoln:mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~ zq ~&�w  bsq ~ '[ac3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�	sq ~ L��Iuq ~ O   q ~q ~ �w  �sq ~ '�8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t miami:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L16�uq ~ O   q ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t charleston:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�'sq ~ L]�uq ~ O   q ~�w  �sq ~ '�]�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~�.q ~�-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�4sq ~ L�O�uq ~ O   q ~<q ~ w  �sq ~ '���0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8=xq ~�;q ~�:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Asq ~ L���uq ~ O   q ~�q ~ �w  �sq ~ 'FS��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~�Hq ~�Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Nsq ~ L3�}�uq ~ O   q ~ Qq ~Uq ~5q ~ �w  �sq ~ 'y�$�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@�xq ~�Uq ~�Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�[sq ~ L1-�uq ~ O   q ~ Qq ~ �q ~q ~#w   osq ~ 'z�a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&Xxq ~�bq ~�asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�hsq ~ L;���uq ~ O   q ~�w  "sq ~ '�E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�oq ~�nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�usq ~ L+
$uq ~ O   q ~ Rq ~ Sq ~ gw  �sq ~ ''q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~o�xq ~�|q ~�{sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L5t�uq ~ O   q ~o�q ~ �w  �sq ~ '�}Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t ohio:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L 4�uq ~ O   q ~�w  �sq ~ '(/,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ixq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�^yuq ~ O   q ~O~w  �sq ~ '� ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���Nuq ~ O   q ~ Qq ~gq ~hw  Isq ~ '.��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~��sq ~ L-��uq ~ O   q ~�w   sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_wilsont mount_wilson:mxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�^v_uq ~ O   q ~ zt wilsonw  �sq ~ '~�%�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"=xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L ��3uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '(~#�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
san_angelot san_angelo:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��L�uq ~ O   q ~ �q ~w  �sq ~ 'H�-Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~IUxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LiU\suq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t newton:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�|3�uq ~ O   q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4�xq ~�	q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�50�uq ~ O   q ~ Qq ~ �q ~$q ~$w  �sq ~ '���>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~2�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�١|uq ~ O   q ~2�w  Xsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~B�t tempe:nxq ~�#q ~�"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�+sq ~ L�7Ouq ~ O   q ~B�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�2q ~�1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~�xq ~�8sq ~ L �uq ~ O   q ~ w   -sq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"�xq ~�?q ~�>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Esq ~ L��0}uq ~ O   q ~
/q ~	�w  sq ~ '�� q ~�sq ~ sq ~ sq ~ J   w   q ~Eq ~5xq ~�Kq ~�Jsq ~ @q ~�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~�Osq ~ L ���uq ~ O   q ~<w  
sq ~ '�׊�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�Vq ~�Usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�\sq ~ L����uq ~ O   q ~ fq ~�w  0sq ~ '�hkxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t troy:nxq ~�cq ~�bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�ksq ~ L 6u&uq ~ O   q ~�w   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~�rq ~�qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�xsq ~ L��ruq ~ O   q ~&�q ~5w  �sq ~ '%���q ~�sq ~ sq ~ sq ~ 
w   q ~Aq ~	!q ~1vxq ~�~q ~�}sq ~ @q ~�sq ~ G)���    sq ~ sq ~ J   w   q ~ �q ~	,q ~ <xq ~��q ~�w   gsq ~ 'zl��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lg�<ouq ~ O   q ~Uq ~5q ~ �w  sq ~ '��Mrsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~P�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lb���uq ~ O   q ~ Rq ~ Sq ~B�w  	,sq ~ 'o�8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~\Pxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L9=�uq ~ O   q ~ Qq ~ �q ~=Ow  ~sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^xxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�J|uq ~ O   q ~Uq ~Ew  sq ~ '<OKMq ~�sq ~ sq ~ sq ~ J   w   q ~Exq ~��q ~��sq ~ @q ~�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~ L��auq ~ O   q ~Ww  
]sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�`G�uq ~ O   q ~�q ~ �w  �sq ~ '�Gysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t great_salt_laket great_salt_lake:lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lc"�uq ~ O   q ~q ~Dq ~q ~w  Osq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t rainyt rainy:lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�˖uq ~ O   q ~q ~��w  �sq ~ '��q ~�sq ~ sq ~ sq ~ J   w   q ~|xq ~��q ~��sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~��sq ~ L 5�@uq ~ O   t spotw  
sq ~ 'cˏ[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�݆Guq ~ O   q ~�q ~�w   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~F.t pittsburgh:nxq ~�
q ~�	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�gj�uq ~ O   q ~F.w  "sq ~ '.��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~o�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L<e�uq ~ O   q ~ Qq ~o�q ~ �w  �sq ~ 'OS;\q ~$�sq ~ sq ~ sq ~ 
w   q ~�xq ~�%q ~�$sq ~ @q ~$�sq ~ G���    sq ~ sq ~ J   w   q ~�xq ~�)q ~%w   Qsq ~ '�w�Esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3�xq ~�.q ~�-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�4sq ~ L�C��uq ~ O   q ~�q ~�q ~Fw  }sq ~ '��9sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5�xq ~�;q ~�:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Asq ~ L_��uq ~ O   q ~Iq ~ Rw  �sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�Hq ~�Gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�Nsq ~ L  �uq ~ O   t byw   sq ~ '�.�jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~�Vq ~�Usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�\sq ~ LE؂uq ~ O   q ~ Qq ~ �q ~'�w  �sq ~ '-f��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~z�xq ~�cq ~�bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�isq ~ L����uq ~ O   q ~?�w  �sq ~ '�nqXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~?t tacoma:nxq ~�pq ~�osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�xsq ~ L�w�+uq ~ O   q ~?w  Tsq ~ 'E"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"�xq ~�q ~�~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L����uq ~ O   q ~ Qq ~"�w  �sq ~ '&�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~1t lynn:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L 2�Kuq ~ O   q ~1w  Psq ~ '  �q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~ L  �uq ~ O   q ~-�w  	�sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t new_britaint new_britain:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L܌+uq ~ O   q ~�q ~tw  �sq ~ '��ոsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�WW�uq ~ O   q ~
�q ~9�q ~ �w  	esq ~ '�\�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~5cxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�9�nuq ~ O   q ~ Qq ~�q ~ �w  �sq ~ 'z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�y�uq ~ O   q ~�w  	�sq ~ 'I�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~f�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L[���uq ~ O   q ~E)q ~w  }sq ~ '�"=bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LL�H�uq ~ O   q ~�q ~B�w  /sq ~ 'E��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�vz�uq ~ O   q ~�q ~Tw  �sq ~ 'yi~�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~04xq ~�q ~� sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L.G%uq ~ O   q ~0?q ~5w   ysq ~ '�w�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L	���uq ~ O   q ~q ~=q ~ �w   �sq ~ '��!�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�!sq ~ Lk��uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ '�ڼ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~<t downey:nxq ~�(q ~�'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�0sq ~ L���uq ~ O   q ~<w   }sq ~ '�"{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~{xq ~�7q ~�6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�=sq ~ Lu�~�uq ~ O   q ~�q ~0�w  sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*oxq ~�Dq ~�Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Jsq ~ L{�Kuq ~ O   q ~*zq ~ �w  "sq ~ '��S�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@�xq ~�Qq ~�Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Wsq ~ L�׾uq ~ O   q ~@�q ~�w  �sq ~ '�̙;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�^q ~�]sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�dsq ~ L���uq ~ O   q ~Xq ~?�w  �sq ~ 'krsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Axq ~�kq ~�jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�qsq ~ LgTPuq ~ O   q ~Lw  #sq ~ '��&�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'xq ~�xq ~�wsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�~sq ~ LzbQ}uq ~ O   q ~2w  �sq ~ 'Y�X�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~6�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�buq ~ O   q ~ Qq ~ �q ~6�w  �sq ~ '�k�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~
�t laredo:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�ץ1uq ~ O   q ~
�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'}t erie:lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LOF�uq ~ O   q ~q ~'}w  Csq ~ '��R�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L@��#uq ~ O   q ~?q ~�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�,S�uq ~ O   q ~�w  �sq ~ 'v��Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�h�tuq ~ O   q ~$�w  nsq ~ 'AI��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	Exq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��+uq ~ O   q ~ Qq ~ �q ~	Pq ~ �w  	gsq ~ '��a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_crestonet mount_crestone:mxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L-�w6uq ~ O   q ~ zq ~EYw  Zsq ~ '��
sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L ��uq ~ O   q ~]w  �sq ~ '�U�jq ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~� q ~��sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�sq ~ LK�ipuq ~ O   t 	traversedw  
(sq ~ '䧽�q ~�sq ~ sq ~ sq ~ J   w   q ~Aq ~Hq ~Hxq ~�q ~�
sq ~ @q ~�sq ~ G���    sq ~ sq ~ J   w   q ~ �q ~q ~xq ~�q ~+$w  	�sq ~ '029Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�7 Auq ~ O   q ~�q ~�q ~5w  "sq ~ '�?J�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^�xq ~�!q ~� sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�'sq ~ Lv�(juq ~ O   q ~ Qq ~^�q ~ �w  	�sq ~ '��q ~W�sq ~ sq ~ sq ~ 
w   q ~Eq ~5xq ~�-q ~�,sq ~ @q ~W�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~�1q ~W�w   1sq ~ '�4�;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-Nxq ~�6q ~�5sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�<sq ~ Lj��uq ~ O   q ~-Yq ~(�w  sq ~ 'Yo�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	lansing:nxq ~�Cq ~�Bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Ksq ~ L���uq ~ O   q ~�w  &sq ~ '��I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<jxq ~�Rq ~�Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Xsq ~ L֍��uq ~ O   q ~ Qq ~ �q ~"Nw  Isq ~ '޺�\sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1�xq ~�_q ~�^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�esq ~ L����uq ~ O   q ~ Qq ~1�q ~ �w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�lq ~�ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�rsq ~ L��22uq ~ O   q ~�q ~�q ~Tw  ksq ~ ';��7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~}xq ~�yq ~�xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Fuq ~ O   q ~�q ~�w  �sq ~ 'h�Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L����uq ~ O   q ~�q ~ �w  sq ~ '�QZ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Dt 
hamilton:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��gzuq ~ O   q ~Dw  �sq ~ '��'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���>uq ~ O   q ~�q ~v�w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�X�uq ~ O   q ~"w  =sq ~ '6]�Vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;;xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�kouq ~ O   q ~;Fq ~w  �sq ~ '@,�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~G�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ La��(uq ~ O   q ~ Qq ~ �q ~�w  9sq ~ 'o�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Vt monroe:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�P'zuq ~ O   q ~Vw  	�sq ~ '�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	!xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~��sq ~ L�Xۇuq ~ O   q ~p�w   
sq ~ '.)JRsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�&�uq ~ O   q ~ Rq ~ Sq ~�w  vsq ~ 't�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~%t flint:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~%w  �sq ~ '�5�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t lower_meriont lower_merion:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L~d$�uq ~ O   q ~)q ~)w  �sq ~ 'ȧWxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~/�t inglewood:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�&sq ~ Ly�Fuq ~ O   q ~/�w  sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)wxq ~�-q ~�,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�3sq ~ Ln���uq ~ O   q ~ Qq ~�q ~�q ~ �w   �sq ~ '�$k{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$6xq ~�:q ~�9sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�@sq ~ L�M�muq ~ O   q ~$Aq ~ �w  isq ~ ' 8#Asq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�Gq ~�Fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�Msq ~ L 7�uq ~ O   t whatw   sq ~ '�jvsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�Uq ~�Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�[sq ~ L�:�uq ~ O   q ~ Qq ~ �q ~�w  |sq ~ 'D	7sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~F#xq ~�bq ~�asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�hsq ~ L;`<uq ~ O   q ~F.q ~w  Jsq ~ '7��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Q�xq ~�oq ~�nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�usq ~ L��uq ~ O   t citiesw   Ksq ~ '��D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t sterling_heightst sterling_heights:nxq ~�}q ~�|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L� ��uq ~ O   q ~�q ~�w  (sq ~ 'F�lq ~�sq ~ sq ~ sq ~ J   w   q ~xq ~��q ~��sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~ L�Z��uq ~ O   t inhabitantsw  
Dsq ~ '�4��q ~�sq ~ sq ~ sq ~ J   w   q ~WRxq ~��q ~��sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~ L 7�uq ~ O   q ~�Pw  	�sq ~ '�FBq ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~ L�E�uq ~ O   t throughw  	�sq ~ 'O��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~f�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lb&�uq ~ O   q ~E)q ~ �w  �sq ~ '�G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t 
beaumont:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LO2�]uq ~ O   q ~w  sq ~ 'W)��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~c#xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��� uq ~ O   q ~c.q ~ �w  �sq ~ '&�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~I�t 
savannah:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�Juq ~ O   q ~I�w   �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L^���uq ~ O   q ~ Qq ~ �q ~�w   �sq ~ '-���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~It 	alabama:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���uq ~ O   q ~Iw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Gt lowell:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��5uq ~ O   q ~Gw  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~f�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��j@uq ~ O   q ~ Qq ~f�q ~g w  �sq ~ 'e(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�!sq ~ L��juq ~ O   q ~�w  �sq ~ '&�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	compton:nxq ~�(q ~�'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�0sq ~ L8��"uq ~ O   q ~�w  
sq ~ '�y@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~�7q ~�6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�=sq ~ Lp��uq ~ O   q ~
w   �sq ~ 'Jt��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	orlando:nxq ~�Dq ~�Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Lsq ~ L�{�uq ~ O   q ~�w  �sq ~ ':�Zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~?�xq ~�Sq ~�Rsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Ysq ~ L.��uq ~ O   q ~ Qq ~ �q ~?�w  jsq ~ '{��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8^xq ~�`q ~�_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�fsq ~ L �-uq ~ O   q ~8iw  *sq ~ '�?]]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~J�xq ~�mq ~�lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�ssq ~ L\>�uq ~ O   q ~
�q ~ �w  ysq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�zq ~�ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���nuq ~ O   q ~�q ~"�w  sq ~ '-�8-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Kxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�!��uq ~ O   q ~Vq ~�w   �sq ~ '1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~5t tennessee:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�@��uq ~ O   q ~5w  �sq ~ '�K!sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LZ
�uq ~ O   q ~�q ~Ew  �sq ~ '[!�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~/t 	clinton:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L3O��uq ~ O   q ~/w  Dsq ~ '�d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	champlaint champlain:lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L[�UJuq ~ O   q ~q ~��w  Ysq ~ '���'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_kennedyt mount_kennedy:mxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�)'�uq ~ O   q ~ zt kennedyw   �sq ~ 'j=�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~)�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�Ruq ~ O   q ~ w  �sq ~ 'K��8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~7�t 	decatur:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L[�Puq ~ O   q ~7�w  �sq ~ '�V��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~M=xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~ Qq ~ �q ~MHw  <sq ~ 'r{Y�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~.Wt 
syracuse:nxq ~�	q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LsOuq ~ O   q ~.Ww  Qsq ~ '�P�[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L 8uq ~ O   q ~ Qq ~]w  qsq ~ 'Ƽ�Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~�%q ~�$sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�+sq ~ LN;��uq ~ O   q ~<q ~"w  Jsq ~ '�L��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~drxq ~�2q ~�1sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�8sq ~ L�)ٓuq ~ O   q ~�q ~ Rw  ]sq ~ 'y�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'t elgin:nxq ~�?q ~�>sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Gsq ~ L��uq ~ O   q ~'w  sq ~ '��kXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~. t evansville:nxq ~�Nq ~�Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Vsq ~ L���uq ~ O   q ~. w  sq ~ '3�Msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�]q ~�\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�csq ~ Lt~%�uq ~ O   q ~�q ~ Rw  �sq ~ '��<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~�jq ~�isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�psq ~ L��uq ~ O   q ~Wq ~"w  {sq ~ '��@�q ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~�vq ~�usq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�zsq ~ LD7�uq ~ O   t 	mountainsw  
Jsq ~ ';��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~4xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��1]uq ~ O   q ~?q ~�w  Rsq ~ 'mLXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ht southfield:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L0,�uq ~ O   q ~Hw  �sq ~ '��_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Uxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�J�uq ~ O   q ~ Qq ~ �q ~ �q ~`w  ^sq ~ 'ʃ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t louisiana:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L~l�uq ~ O   q ~�w  �sq ~ '-
�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#0xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��ۭuq ~ O   q ~�q ~ �w  sq ~ '�9Fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!exq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��{wuq ~ O   q ~�w  �sq ~ '��]^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	Vxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LRy�Buq ~ O   q ~ Qq ~ �q ~	aq ~	bw  sq ~ '��R_sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��Wuq ~ O   q ~�w   �sq ~ '�y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t connecticut:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lf�1auq ~ O   q ~�w  0sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~cxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LA��Kuq ~ O   q ~nq ~w  �sq ~ 'G.�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t salt_lake_cityt salt_lake_city:nxq ~�
q ~�	sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~q ~q ~ �w  |sq ~ ')��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~G#xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~� sq ~ L��~�uq ~ O   q ~G.q ~w  6sq ~ '���wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�'q ~�&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�-sq ~ L3L�uq ~ O   q ~�w  	rsq ~ 'pX�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�4q ~�3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�:sq ~ LV���uq ~ O   q ~�q ~�w  Xsq ~ 'r��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~}xq ~�Aq ~�@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Gsq ~ L�9�uq ~ O   q ~�q ~Tw  �sq ~ '`-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~>t middletown:nxq ~�Nq ~�Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Vsq ~ L�Lq�uq ~ O   q ~>w  sq ~ 'a�<sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~�]q ~�\sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�csq ~ L�D�uq ~ O   q ~ Qq ~q ~ �w  �sq ~ '��s�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~�jq ~�isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�psq ~ L�z��uq ~ O   q ~Mq ~ Rw  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
�xq ~�wq ~�vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�}sq ~ L�B��uq ~ O   q ~
�w  sq ~ 't; >sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��uq ~ O   q ~+w  Ysq ~ '�N�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t sunnyvale:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�*#9uq ~ O   q ~�w  Esq ~ '�ؚ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~*oxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L����uq ~ O   q ~ Qq ~ �q ~*zw  Msq ~ '<,��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�l��uq ~ O   q ~ Qq ~ �q ~�w  �sq ~ 'Q�csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~fxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L`��uq ~ O   q ~ Qq ~ Rq ~ Sq ~gw  +sq ~ '��tq ~�sq ~ sq ~ sq ~ J   w   q ~Mxq ~��q ~��sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~ L 7�uq ~ O   q ~w  
Wsq ~ 'w�h�q ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~��q ~��sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~ L  �uq ~ O   q ~jw  
Isq ~ '��ƙsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~dxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�d�uq ~ O   q ~ Qq ~Nq ~d&w  	�sq ~ 'Qo/sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�K)�uq ~ O   q ~q ~ �q ~�w  
sq ~ 'Orsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L훈uq ~ O   q ~ Qq ~ �q ~ q ~;w  |sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~@�t largo:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�
sq ~ L��uq ~ O   q ~@�w  �sq ~ 'n�B�q ~O�sq ~ sq ~ sq ~ 
w   q ~Exq ~�q ~�sq ~ @q ~O�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~�q ~O�w   sq ~ 'k�esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A"xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�y>�uq ~ O   q ~A-w  zsq ~ '�
�osq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~pxq ~�&q ~�%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�,sq ~ L~�lXuq ~ O   q ~{w  �sq ~ '� ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~�3q ~�2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�9sq ~ L  huq ~ O   q ~z�w   3sq ~ '�B�Ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~�@q ~�?sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Fsq ~ L�g��uq ~ O   q ~)w  	�sq ~ '�2��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.�xq ~�Mq ~�Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Ssq ~ L��Njuq ~ O   q ~.�q ~w  %sq ~ '1*sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�Zq ~�Ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�`sq ~ L=xf}uq ~ O   q ~ Qq ~ �q ~ �w   �sq ~ '�)_�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t irvington:nxq ~�gq ~�fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�osq ~ L-�Yuq ~ O   q ~w  sq ~ 'F���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~pAxq ~�vq ~�usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�|sq ~ L�UNTuq ~ O   q ~ �q ~CCq ~ �w   �sq ~ 'w<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�y�uq ~ O   q ~Nq ~�q ~w  �sq ~ '_l�Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��t[uq ~ O   q ~�q ~!q ~�w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LϢ!uq ~ O   q ~yq ~"w  sq ~ ' 3)q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~ L 2��uq ~ O   t listw  
:sq ~ '5���q ~�sq ~ sq ~ sq ~ J   w   q ~Eq ~Hxq ~��q ~��sq ~ @q ~�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~��sq ~ L��y�uq ~ O   t tallestw  
	sq ~ 'V��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~h@xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L*
�uq ~ O   q ~q ~Cq ~�w  ?sq ~ '0p�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�-��uq ~ O   q ~ Rq ~ Sq ~q ~ w  Esq ~ '~hϘsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~(�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��uq ~ O   q ~
�q ~(�q ~w  sq ~ '*¼sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L k��uq ~ O   q ~ Qq ~�w  �sq ~ 'Ttv�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LT��uq ~ O   q ~�q ~ �w  �sq ~ 'w��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LK��auq ~ O   q ~Fq ~ �w  �sq ~ 'bO�isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~q ~�q ~Fw  *sq ~ 'ŜBssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�P%uq ~ O   q ~ >q ~ Rw  nsq ~ '�'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_shavanot mount_shavano:mxq ~�&q ~�%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�/sq ~ L:��?uq ~ O   q ~ zt shavanow  �sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~�7q ~�6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�=sq ~ LE��uq ~ O   q ~ Rq ~ Sq ~w  qsq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~AKt 
metairie:nxq ~�Dq ~�Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Lsq ~ L�/��uq ~ O   q ~AKw  �sq ~ ' 1�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~�Tsq ~ L �Vuq ~ O   q ~�w  
sq ~ '�l�msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~#hxq ~�[q ~�Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�asq ~ L�S�fuq ~ O   q ~#sq ~ �w  �sq ~ '��esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�hq ~�gsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�nsq ~ L�4uq ~ O   q ~ Qq ~ �q ~�w  wsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!Ixq ~�uq ~�tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�{sq ~ L����uq ~ O   q ~fw  �sq ~ '4��usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��p�uq ~ O   q ~�q ~ Rw  �sq ~ '�U�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LC{ٓuq ~ O   q ~
q ~ �w  �sq ~ '��bsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��uq ~ O   q ~ Qq ~ �q ~ww  �sq ~ '� @sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�Vuq ~ O   q ~ fq ~�q ~ gw  	4sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lb�uq ~ O   q ~ �q ~9�w  	6sq ~ '?�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~%�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L5o�uq ~ O   q ~q ~q ~"w  sq ~ '���~sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Rxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Li�uq ~ O   q ~ Qq ~ �q ~]q ~	w  	7sq ~ '�3�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~>�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�? uq ~ O   q ~ Qq ~>�q ~ �w  ^sq ~ '�?�wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L����uq ~ O   q ~�w  7sq ~ 'POr�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~E�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~ L�~�Cuq ~ O   q ~o�w   "sq ~ 'X&�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�
sq ~ L^�@uq ~ O   q ~ Qq ~ �q ~gq ~/q ~0w  %sq ~ 'i{#8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Lt huntsville:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LgTPuq ~ O   q ~Lw  	sq ~ '�O�Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~$�xq ~� q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�&sq ~ L��*uq ~ O   q ~hq ~"w  rsq ~ '"��xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 
stamford:nxq ~�-q ~�,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�5sq ~ LN0$�uq ~ O   q ~�w  8sq ~ '���[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,�xq ~�<q ~�;sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Bsq ~ L��uq ~ O   q ~,�q ~pw  �sq ~ '�rBAsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~�Iq ~�Hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Osq ~ L���uq ~ O   q ~q ~=q ~	bq ~�w  �sq ~ '�,َsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�Vq ~�Usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�\sq ~ LC�8uq ~ O   q ~ Qq ~ �q ~q ~ �w   sq ~ ':��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~h@xq ~�cq ~�bsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�isq ~ L�pGuq ~ O   q ~q ~Cw  	@sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ 4xq ~�pq ~�osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�vsq ~ L���uq ~ O   q ~ Rq ~ Sq ~ >w  Vsq ~ ' )�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~�~sq ~ L �[uq ~ O   t perw  	�sq ~ 'Kłsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!Ixq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L>Å�uq ~ O   q ~fq ~ Rw  lsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LN�Z�uq ~ O   q ~ Qq ~ �q ~�q ~�w  Asq ~ '//�Vsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&ixq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L,b�yuq ~ O   q ~ Qq ~ �q ~�q ~ �w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~'Jt 	memphis:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L8�0�uq ~ O   q ~'Jw   �sq ~ 'g���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&ixq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Ld�~�uq ~ O   q ~�q ~ �q ~�w  �sq ~ 'zG�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~{xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L?C�uq ~ O   q ~�q ~5w   �sq ~ '��SUsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�uuq ~ O   q ~�q ~�q ~�w  Rsq ~ ' 3�q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~ L 3z�uq ~ O   t namew  	�sq ~ '���+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t naknekt naknek:lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�]�uq ~ O   q ~q ~��w  Hsq ~ 'B��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Eq ~	!xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~�sq ~ L i�uq ~ O   q ~ Qq ~w   Zsq ~ 'ڗR5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~�	q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��uq ~ O   q ~q ~"w  8sq ~ '�&�+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�F6uq ~ O   q ~�q ~�w  Esq ~ '��6�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�#q ~�"sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�)sq ~ L��6 uq ~ O   q ~Xw  	Osq ~ 'm�c�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~@+xq ~�0q ~�/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�6sq ~ L��1Juq ~ O   q ~�q ~�w  lsq ~ 'yUsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 	santa_anat santa_ana:nxq ~�=q ~�<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Fsq ~ L��uuq ~ O   q ~ q ~$w  ^sq ~ '�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Mt district_of_columbia:nxq ~�Mq ~�Lsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Usq ~ L���wuq ~ O   q ~Wq ~ Sq ~Xw  �sq ~ '֒;�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Uxq ~�\q ~�[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�bsq ~ L��'@uq ~ O   q ~ �q ~`q ~"w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�iq ~�hsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�osq ~ L\=uq ~ O   q ~ Qq ~�q ~�q ~ �w  >sq ~ 'y���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ Nt salem:nxq ~�vq ~�usq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�~sq ~ L�IDuq ~ O   q ~ Nw  tsq ~ '�"9Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�F�uq ~ O   q ~�q ~ �w  �sq ~ 'R���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LYDxuq ~ O   q ~ �q ~ �w  �sq ~ ',b��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~+�t 
scranton:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�C3buq ~ O   q ~+�w  sq ~ 'F�'sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ut akron:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�E�uq ~ O   q ~uw  �sq ~ '0	�wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t st_louist 
st_louis:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L'�uq ~ O   q ~Nq ~w  )sq ~ '3BY�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~;xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�jO�uq ~ O   q ~ Qq ~ �q ~Fw  	sq ~ 'o�|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~]xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lh�Euq ~ O   q ~ Qq ~ �q ~hw  �sq ~ ')y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���uq ~ O   q ~<w  �sq ~ '�(sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~yt fullerton:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�^��uq ~ O   q ~yw  Xsq ~ '�TX�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�	sq ~ L �uq ~ O   q ~ Qq ~�q ~�w  sq ~ '@u�`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lr�c�uq ~ O   q ~ Qq ~ �q ~�w  &sq ~ 'Hbsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A@xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�#sq ~ L��uq ~ O   q ~AKq ~"�w   �sq ~ 'P{2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~<Lxq ~�*q ~�)sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�0sq ~ L��v�uq ~ O   q ~ Rq ~ Sq ~3w  ^sq ~ 'ԩ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�7q ~�6sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�=sq ~ L���uq ~ O   q ~�w  �sq ~ '�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~I�xq ~�Dq ~�Csq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Jsq ~ L�Juq ~ O   q ~I�w  Osq ~ '�)'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~qt 
richmond:nxq ~�Qq ~�Psq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Ysq ~ L����uq ~ O   q ~qw  �sq ~ '�V�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t miami_beacht miami_beach:nxq ~�`q ~�_sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�isq ~ LŊ�uq ~ O   q ~�q ~	bw  _sq ~ 'dt�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"exq ~�pq ~�osq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�vsq ~ L��3uq ~ O   q ~?w  _sq ~ '�ZXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~�}q ~�|sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���wuq ~ O   q ~Wq ~ Sq ~Xw  @sq ~ '�/m�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~pxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L;�!�uq ~ O   q ~{q ~"w  qsq ~ '% �q ~�sq ~ q ~Swq ~Swsq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��q ~�w  
sq ~ '��0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���uq ~ O   q ~3q ~'�q ~=w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t 	hampton:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L)Bӵuq ~ O   q ~�w  -sq ~ 'ȣ�0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LC�uq ~ O   q ~Wq ~ �w  Nsq ~ '>�iZsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��Tuq ~ O   q ~ �q ~�q ~ �w  �sq ~ '��m[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Jxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�"8Euq ~ O   q ~Uq ~	�w  �sq ~ '��6,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~J�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lb��uq ~ O   q ~ Qq ~
�q ~ �w  Lsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~1�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�|uq ~ O   q ~ �q ~1�q ~w  Csq ~ '��a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~drxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~� sq ~ L^��uq ~ O   q ~ Qq ~ Rq ~ Sq ~�w  �sq ~ '�Օ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~Uw   wsq ~ 'aDuysq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~vxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LFLG�uq ~ O   q ~�w  sq ~ 'tV8xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~.�t bethlehem:nxq ~�!q ~� sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�)sq ~ Lm�s�uq ~ O   q ~.�w  �sq ~ '�1C�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~"xq ~�0q ~�/sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�6sq ~ L|�+(uq ~ O   q ~#q ~ Rw  Qsq ~ 'K�q ~�sq ~ sq ~ sq ~ J   w   sq ~ 0q ~ :t death_valleyt death_valley:loxq ~�<q ~�;sq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Csq ~ L��{�uq ~ O   q ~w  
sq ~ 'E�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~{t 	norwalk:nxq ~�Jq ~�Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Rsq ~ L~�lXuq ~ O   q ~{w  �sq ~ '��O�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[Lxq ~�Yq ~�Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�_sq ~ LO6�uq ~ O   q ~[Ww  bsq ~ '�T��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~t 	altoona:nxq ~�fq ~�esq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�nsq ~ L���uq ~ O   q ~w   �sq ~ 'և[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~�uq ~�tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�{sq ~ L���uq ~ O   q ~�q ~Fw  �sq ~ 'M7�5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�&nuq ~ O   q ~ Qq ~ �q ~!�w  �sq ~ '
�O�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�2\�uq ~ O   q ~�q ~=w  #sq ~ '%�/sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~J}xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L �vZuq ~ O   q ~gw  �sq ~ '�`=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LR`6suq ~ O   q ~�w  qsq ~ 'd��q ~]sq ~ sq ~ sq ~ 
w   q ~�q ~Hxq ~��q ~��sq ~ @q ~]sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~��q ~]w   Tsq ~ '<��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��uq ~ O   q ~ Qq ~ �q ~�w  asq ~ 'Ɯ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lr��uq ~ O   q ~ Qq ~ �q ~�w  ,sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L6.�luq ~ O   q ~ Rq ~ Sq ~5w  `sq ~ '�G�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~'Pxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L5y�uq ~ O   q ~ Qq ~ �q ~'[w  �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ Lž�uq ~ O   q ~-�w  Isq ~ '5�f�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��4�uq ~ O   q ~ Qq ~ �q ~&w  fsq ~ '�}��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L����uq ~ O   q ~ Qq ~ Rq ~ Sq ~�q ~�w  ,sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L1�+uq ~ O   q ~q ~ Rw   �sq ~ '��x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~z�xq ~�&q ~�%sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�,sq ~ L�9`�uq ~ O   q ~?�q ~ �w  �sq ~ '��kUsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^xxq ~�3q ~�2sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�9sq ~ LJ���uq ~ O   q ~ Qq ~ �q ~Uq ~Ew  �sq ~ '=�Nq ~�sq ~ sq ~ sq ~ J   w   q ~�xq ~�?q ~�>sq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�Csq ~ L 6M�uq ~ O   q ~*w  
`sq ~ '�p�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�Jq ~�Isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Psq ~ L�n�uq ~ O   q ~ Rq ~ Sq ~�w  Dsq ~ '��S�q ~�sq ~ sq ~ sq ~ J   w   q ~Q�xq ~�Vq ~�Usq ~ @q ~�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~�Zsq ~ L   �uq ~ O   q ~�w  
Fsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Sxq ~�aq ~�`sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�gsq ~ Lx��8uq ~ O   q ~^q ~Uq ~�w  �sq ~ 'VR{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�nq ~�msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�tsq ~ L�փ�uq ~ O   q ~ �q ~�q ~iw  9sq ~ '�F]�q ~�sq ~ sq ~ sq ~ J   w   q ~xq ~�zq ~�ysq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~�~sq ~ L���uq ~ O   q ~ Rw  
.sq ~ '2�^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~ L�b�uq ~ O   q ~w   \sq ~ '��^�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~	hxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L f�3uq ~ O   q ~�q ~	sw  zsq ~ 'ǫ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~/yxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�[�6uq ~ O   q ~/�q ~ �w  7sq ~ '��q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��q ~uw  	�sq ~ 'y'�Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~&�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�L<uq ~ O   q ~ Qq ~ �q ~&�q ~�w  %sq ~ 'y�Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~!�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�.X�uq ~ O   q ~!�q ~w  �sq ~ '��%sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Zxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L  �uq ~ O   q ~hw  csq ~ '��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~bxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L7��]uq ~ O   q ~Kq ~"�w  csq ~ 'a��[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t cherry_hillt cherry_hill:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L,v��uq ~ O   q ~&�q ~�w  �sq ~ 'q'�"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���&uq ~ O   q ~ Qq ~ �q ~�q ~�w  sq ~ '�D�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�	sq ~ L���"uq ~ O   q ~ Qq ~ �q ~�q ~�w  	Nsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7�xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�5�uq ~ O   q ~7�q ~Uw  Psq ~ '}X�xq ~�sq ~ sq ~ sq ~ J   w   q ~ �xq ~�q ~�sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~� sq ~ L��~uq ~ O   t crossw  
7sq ~ '\�{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�(q ~�'sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�.sq ~ L]t�1uq ~ O   q ~ Qq ~ �q ~
Yw   �sq ~ '�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~afxq ~�5q ~�4sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�;sq ~ L�3�uq ~ O   q ~ Rq ~ Sq ~}w  �sq ~ 'mjP3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
$xq ~�Bq ~�Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Hsq ~ L����uq ~ O   q ~
/w  �sq ~ 'aH&�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~A"xq ~�Oq ~�Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Usq ~ L®�)uq ~ O   q ~A-q ~ �w  �sq ~ 'S<2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~7 xq ~�\q ~�[sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�bsq ~ L`\�uq ~ O   q ~�t dcw  �sq ~ '9sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t new_orleanst new_orleans:nxq ~�jq ~�isq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�ssq ~ L��
uq ~ O   q ~�q ~!w  �sq ~ 'eDl�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.Lxq ~�zq ~�ysq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L���uq ~ O   q ~.Wq ~�w  �sq ~ ' 6�.q ~�sq ~ q ~�q ~�sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~ L 6C�uq ~ O   q ~-�w  	�sq ~ 'ܑ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�OPuq ~ O   q ~ �q ~q ~w  �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Ft springfield:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�1�Kuq ~ O   q ~Fw  	msq ~ 'Qq�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~-�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��5�uq ~ O   q ~ Qq ~ �q ~. w  �sq ~ '&[e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L��E�uq ~ O   q ~ �q ~�q ~Aw  �sq ~ '���;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t port_arthurt port_arthur:nxq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L�aWAuq ~ O   q ~!�q ~!�w  2sq ~ '3"��q ~�sq ~ sq ~ sq ~ J   w   q ~Hxq ~��q ~��sq ~ @q ~�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~ L 0��uq ~ O   q ~�w  	�sq ~ 'Ǳ0sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ixq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ L����uq ~ O   q ~O~q ~ �w  6sq ~ '�B��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~0	xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LV�vuq ~ O   q ~0w  �sq ~ '��=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~><xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~��sq ~ LAֳ�uq ~ O   q ~ Qq ~ �q ~*w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t 
south_bendt south_bend:nxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lʾ��uq ~ O   q ~
�q ~(�w  �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ nt mount_grayst mount_grays:mxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�4Wuq ~ O   q ~ zt graysw  isq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~dxq ~�'q ~�&sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�-sq ~ LN��uq ~ O   q ~oq ~pq ~w  	�sq ~ '��;sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~L�xq ~�4q ~�3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�:sq ~ L�uXuq ~ O   q ~B�q ~w  sq ~ '^�Gsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~bjxq ~�Aq ~�@sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Gsq ~ L�W�Suq ~ O   q ~buq ~ �w  �sq ~ '~��Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~=xq ~�Nq ~�Msq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�Tsq ~ L��&uq ~ O   q ~q ~=q ~	bq ~"w  �sq ~ 'WM�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~3�xq ~�[q ~�Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�asq ~ L���uq ~ O   q ~3�q ~pq ~ �w  �xsq ~ !        sq ~ #    ?@      xsq ~ #    ?@     Usr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.LexicalTemplateg��%��	 I hashCodeL 	argumentsq ~ L 
propertiesq ~ (L 	signatureq ~ )L templatet 0Ledu/cornell/cs/nlp/spf/ccg/categories/Category;xpw%�bsq ~ sq ~ sq ~ 
w    xq ~�lq ~�ksq ~ @q ~�Jsq ~ G  �    sq ~ sq ~ J    w    xq ~�psr 5edu.cornell.cs.nlp.spf.ccg.categories.ComplexCategory�f�Ք�nl I hashCodeCacheL syntaxt <Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/ComplexSyntax;xr .edu.cornell.cs.nlp.spf.ccg.categories.CategorycK=�.A� L 	semanticst Ljava/lang/Object;xpsr 'edu.cornell.cs.nlp.spf.mr.lambda.Lambda��Kβ�� L argumentt +Ledu/cornell/cs/nlp/spf/mr/lambda/Variable;L bodyt 4Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L typet 5Ledu/cornell/cs/nlp/spf/mr/language/type/ComplexType;xq ~ 3sr )edu.cornell.cs.nlp.spf.mr.lambda.Variable�u#$rP L 	singletonq ~ xq ~ 1q ~sr 5it.unimi.dsi.fastutil.objects.ReferenceSets$Singleton�7y�J| L elementq ~�txpq ~�|sq ~�vsq ~�{q ~ <sq ~�}q ~��sr (edu.cornell.cs.nlp.spf.mr.lambda.Literalŕtb��� [ 	argumentst 5[Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L 	predicateq ~�x[ 	signaturet /[Ledu/cornell/cs/nlp/spf/mr/language/type/Type;L typeq ~ 2xq ~ 3ur 5[Ledu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression;|�㰢�[i  xp   q ~��sr ;it.unimi.dsi.fastutil.objects.ReferenceSets$UnmodifiableSet�7y�J|  xr Iit.unimi.dsi.fastutil.objects.ReferenceCollections$UnmodifiableCollection�7y�J| L 
collectiont 3Lit/unimi/dsi/fastutil/objects/ReferenceCollection;xpsr 2it.unimi.dsi.fastutil.objects.ReferenceOpenHashSet         F fI sizexp?@     q ~��q ~�|xq ~�|ur /[Ledu.cornell.cs.nlp.spf.mr.language.type.Type;>L5��  xp   q ~ <q ~ <sq ~��sq ~��?@     q ~�|xq ~sr 4it.unimi.dsi.fastutil.objects.ReferenceSets$EmptySet�7y�J|  xpsq ~ ��T��t <<e,e>,<e,e>>q ~q ~w%��sr :edu.cornell.cs.nlp.spf.ccg.categories.syntax.ComplexSyntax$���q\P^ I hashCodeI 	numSlahesL leftt 5Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax;L rightq ~��L slasht 4Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Slash;xr 3edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntaxʊ�	�|��  xp�z�M   sr @edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntax$SimpleSyntax��eBg� I hashCodeL 	attributeq ~ L labelq ~ xq ~�� 3�kt nonet Nq ~��sr 2edu.cornell.cs.nlp.spf.ccg.categories.syntax.Slashѕ�����> C cxp /w   'sq ~�gIH�xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t #0<e,t>t #0<e,t>:<e,t>xq ~��q ~��sq ~ @q ~��sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��q ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��xsq ~ 0sr <edu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType&��M
� I minArgsZ orderSensitiveL optiont ELedu/cornell/cs/nlp/spf/mr/language/type/RecursiveComplexType$Option;xq ~ �l�6�t <t*,t>q ~ �q ~ �    sr Cedu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType$Option�^g� �� Z isOrderSensitiveI 
minNumArgsxp    q ~^t 
and:<t*,t>uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��sq ~ �JW`Lt <<e,t>,<e,t>>q ~ �q ~ �R:L]sq ~���z�M   q ~��q ~��q ~��w   Dsq ~�g 	��sq ~ sq ~ sq ~ 
w   sq ~ 0q ~Tt #0<<e,t>,<<e,e>,e>>t %#0<<e,t>,<<e,e>,e>>:<<e,t>,<<e,e>,e>>xq ~��q ~��sq ~ @q ~nsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vsq ~�{q ~Jsq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~5uq ~��   q ~ :q ~q ~��q ~Jq ~��q ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��xq ~	,q ~��sq ~ �q~Et <<e,t>,<<e,t>,e>>q ~ �q ~	,sq ~��sq ~��?@      xsq ~ �˹�)t <<e,i>,<<e,t>,<<e,t>,e>>>q ~Jq ~����Esq ~���]�   sq ~���ƥY   sq ~�� 4�wq ~��t NPq ~��q ~��sq ~�� 4��q ~��t PPq ~��w   *sq ~�g�K�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t #0<e,<e,t>>t #0<e,<e,t>>:<e,<e,t>>sq ~ 0q ~t #0<e,e>t #0<e,e>:<e,e>sq ~ 0q ~t #1<e,e>t #1<e,e>:<e,e>xq ~�q ~�sq ~ @q ~Lsq ~ G���    sq ~ sq ~ J   w   q ~ �q ~q ~xq ~�sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~� sq ~�vsq ~�{q ~ <sq ~�}q ~�#sq ~��uq ~��   sq ~��uq ~��   q ~�#q ~�$q ~�uq ~��   q ~ <q ~ <sq ~��uq ~��   q ~� q ~�!q ~�uq ~��   q ~ <q ~ <sq ~��sq ~��?@     q ~�#q ~� xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ �$��sq ~���P�   q ~�q ~�	q ~��w   @sq ~�g���sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ <t #0et #0e:exq ~�6q ~�5sq ~ @q ~ �sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�=sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�@sq ~�vsq ~�{q ~ <sq ~�}q ~�Csq ~��uq ~��   sq ~��uq ~��   q ~�Cq ~�7q ~�Dq ~ �uq ~��   q ~ :q ~ :q ~ �sq ~��uq ~��   q ~�Csq ~��sq ~��?@     q ~�Cq ~�@xq ~�@uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�Cq ~�@xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�@xq ~ �q ~��q ~��s-HUsq ~���z�M   q ~��q ~��q ~��w   =sq ~�g�2.dsq ~ sq ~ sq ~ 
w   q ~��xq ~�Xq ~�Wsq ~ @q ~�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~�\sq ~�qsq ~�vsq ~�{q ~sq ~�}q ~�_sq ~�vsq ~�{q ~ �sq ~�}q ~�bsq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�gsq ~��uq ~��   q ~�gsq ~��sq ~��?@     q ~�gq ~�bxq ~�buq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�bxq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~�qsq ~��uq ~��   q ~�qsq ~��sq ~��?@     q ~�_q ~�qxq ~�_uq ~��   q ~ <q ~ <sq ~��sq ~��?@     q ~�_xq ~sq ~��sq ~��?@     q ~�_q ~�bxq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~�_xq ~	,q ~��sq ~ �wй�t <<e,e>,<<e,t>,e>>q ~q ~	,!���sq ~������   sq ~���ƥY   q ~�	q ~��q ~��q ~��q ~��w   sq ~�g�уsq ~ sq ~ sq ~ 
w   q ~�q ~�7xq ~��q ~��sq ~ @q ~�sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��xq ~ �q ~��q ~	!uq ~��   q ~ �q ~q ~�7q ~��q ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xsq ~ ����t <<e,<e,t>>,<e,t>>q ~ �q ~ �q ~��sq ~ ��"(tt <<e,t>,<<e,<e,t>>,<e,t>>>q ~ �q ~��.r�sq ~���7F   sq ~����   sq ~��ȠU�   sq ~�� 3�q ~��t Sq ~�	sq ~�� \sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��q ~��q ~��q ~��w   7sq ~�g���5sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @q ~^^sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��q ~��q ~��q ~��}Usq ~���|�   q ~��q ~��q ~��w   &sq ~�g~��sq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @q ~-sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��xq ~ �q ~�q ~	!uq ~��   q ~ �q ~sq ~��sq ~��?@     q ~��q ~��xq ~Jsq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~	,sq ~��sq ~��?@     q ~��xsq ~ ��Ї�t <<e,<e,t>>,<<e,t>,e>>q ~ �q ~	,q ~��sq ~ �{�t <<e,t>,<<e,<e,t>>,<<e,t>,e>>>q ~ �q ~��8sq ~���<�   sq ~����;!   sq ~���ƥ�   q ~�	q ~��q ~��sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��q ~��q ~��q ~��w   sq ~�g�գ�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�"sq ~�vsq ~�{q ~ <sq ~�}q ~�%sq ~��uq ~��   q ~�%sq ~��sq ~��?@     q ~�%q ~�"xq ~�"uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�"xq ~ �q ~��q ~���՟�sq ~��mLߍ   sq ~��ȠU�   q ~��q ~�	q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��w   sq ~�g<��sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~�4q ~�3sq ~ @q ~Lsq ~ Go��    sq ~ sq ~ J   w   q ~q ~xq ~�8sq ~�qsq ~�vq ~� sq ~�vq ~�#sq ~��uq ~��   sq ~��uq ~��   q ~�#q ~�$q ~�uq ~��   q ~ <q ~ <sq ~��uq ~��   q ~� q ~�!q ~�uq ~��   q ~ <q ~ <sq ~��sq ~��?@     q ~�#q ~� xq ~Auq ~��   q ~q ~q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ �BEq ~�2w   0sq ~�g&���sq ~ sq ~ sq ~ 
w    xq ~�Lq ~�Ksq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�Rsq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�Usq ~�vsq ~�{q ~ �sq ~�}q ~�Xsq ~�vsq ~�{q ~ <sq ~�}q ~�[sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�`sq ~��uq ~��   sq ~��uq ~��   q ~�`sq ~��sq ~��?@     q ~�Uq ~�`xq ~�Uuq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�`q ~�[sq ~��sq ~��?@     q ~�[q ~�Xq ~�`xq ~�Xuq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~�Uq ~�[q ~�Xq ~�`xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�[q ~�Uq ~�Xxq ~ �q ~�qsq ~ 0sq ~ �I:�et 	<<e,t>,t>q ~ �q ~ �t existst exists:<<e,t>,t>uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~�Xq ~�Uxq ~ �sq ~��sq ~��?@     q ~�Uxq ~��q ~��q ~��&���sq ~��x�X�   sq ~���&,�   q ~��sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��q ~��q ~��q ~��w   sq ~�gȨ�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~�uq ~��   q ~ �q ~Jq ~ <q ~��q ~	,��9�sq ~���ƥY   q ~�	q ~��q ~��w   Csq ~�giQsq ~ sq ~ sq ~ 
w   q ~�sq ~ 0q ~	,t #0<<e,t>,e>t #0<<e,t>,e>:<<e,t>,e>xq ~��q ~��sq ~ @q ~�sq ~ G�ǂ    sq ~ sq ~ J   w   q ~ �q ~	,xq ~��sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��q ~��uq ~��   q ~ �q ~ <q ~1vq ~��q ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~��hIqq ~��w   Msq ~�g��{@sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~s~sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~ ��9��sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��w   sq ~�g��{@sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~hosq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~ ��9��sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��w   sq ~�g(�sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @q ~F
sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~��(�>sq ~���|��   q ~��q ~��q ~��w   sq ~�gx�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�
sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�sq ~��uq ~��   q ~�sq ~��sq ~��?@     q ~�q ~�xq ~�uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�xq ~ �q ~�sq ~ 0q ~	,q ~ Qt the:<<e,t>,e>uq ~��   q ~ �q ~ <q ~��q ~	,x~'sq ~���ƥY   q ~�	q ~��q ~��w    sq ~�g(�Ysq ~ sq ~ sq ~ 
w    xq ~�"q ~�!sq ~ @q ~nFsq ~ G  �    sq ~ sq ~ J    w    xq ~�&sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�)sq ~�vsq ~�{q ~ <sq ~�}q ~�,sq ~��uq ~��   q ~�,sq ~��sq ~��?@     q ~�)q ~�,xq ~�)uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�)xq ~ �q ~��q ~��(�ysq ~���|�(   q ~��q ~��q ~��w   sq ~�gV�$�sq ~ sq ~ sq ~ 
w   q ~��xq ~�9q ~�8sq ~ @q ~]sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~�=sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�@sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�Esq ~��uq ~��   q ~�Esq ~��sq ~��?@     q ~�Eq ~�@xq ~�@uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�@xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~�Osq ~��uq ~��   q ~�Oq ~�Pq ~Huq ~��   q ~ :q ~q ~��q ~Jq ~�Lq ~��uq ~��   q ~ �q ~q ~ <q ~��q ~	,�j�sq ~���ƥY   q ~�	q ~��q ~��w   -sq ~�g�y��sq ~ sq ~ sq ~ 
w   q ~��xq ~�Yq ~�Xsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~�_sq ~�qsq ~�vsq ~�{q ~sq ~�}q ~�bsq ~�vsq ~�{q ~ �sq ~�}q ~�esq ~�vsq ~�{q ~ �sq ~�}q ~�hsq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�msq ~��uq ~��   sq ~��uq ~��   q ~�msq ~��sq ~��?@     q ~�eq ~�mxq ~�euq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�msq ~��sq ~��?@     q ~�mq ~�hxq ~�huq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�eq ~�mq ~�hxq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�eq ~�hxq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~�bxq ~�buq ~��   q ~ <q ~ <sq ~��sq ~��?@     q ~�bxq ~sq ~��sq ~��?@     q ~�eq ~�bq ~�hxq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~�eq ~�bxq ~	,sq ~��sq ~��?@     q ~�bxq ~�q ~��sq ~ ��U�%t <<e,e>,<<e,t>,<<e,t>,e>>>q ~q ~�\�sq ~��(��O   sq ~���]�   sq ~���ƥY   q ~�	q ~��q ~��q ~�q ~��q ~��q ~��w   ,sq ~�gEH=sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~ �D�t�sq ~��ȠU�   q ~��q ~�	q ~��w   )sq ~�g�q��sq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��q ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~�ʗc$�sq ~���k�   q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��w   <sq ~�gI�Gmsq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @q ~��sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ <sq ~��sq ~��?@     q ~��xq ~sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��xq ~Vq ~��q ~T�a��sq ~������   sq ~���ƥ�   q ~�	q ~��q ~��q ~��q ~��w   sq ~�g䤶�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~-sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~�sr 4edu.cornell.cs.nlp.spf.ccg.categories.SimpleCategory��4_C� I hashCodeCacheL syntaxt BLedu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax$SimpleSyntax;xq ~�ssq ~�vsq ~�{q ~ <sq ~�}q ~�sq ~��uq ~��   q ~�q ~�q ~�uq ~��   q ~ <q ~ <q ~��q ~���yq ~��w   6sq ~�g�;�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�sq ~�vsq ~�{q ~ �sq ~�}q ~�sq ~�vsq ~�{q ~ <sq ~�}q ~�sq ~��uq ~��   sq ~��uq ~��   q ~�sq ~��sq ~��?@     q ~�q ~�xq ~�uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�sq ~��sq ~��?@     q ~�q ~�xq ~�uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�q ~�q ~�xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�q ~�xq ~ �sq ~��sq ~��?@     q ~�xq ~��q ~��sq ~ �˪xt <<e,t>,<<e,t>,<e,t>>>q ~ �q ~�ʕ;�%sq ~��8���   sq ~���f   q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��q ~��q ~��w   3sq ~�gGsJ�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t #0<t,t>t #0<t,t>:<t,t>xq ~�;q ~�:sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G���    sq ~ sq ~ J   w   q ~�xq ~�Dsq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�Gsq ~�vsq ~�{q ~ <sq ~�}q ~�Jsq ~��uq ~��   sq ~��uq ~��   q ~�Jsq ~��sq ~��?@     q ~�Jq ~�Gxq ~�Guq ~��   q ~ <q ~ �q ~�Pq ~�<uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~�Gxq ~ �q ~��q ~��|�[�sq ~���z�M   q ~��q ~��q ~��w   ?sq ~�g:��sq ~ sq ~ sq ~ 
w   q ~��xq ~�Zq ~�Ysq ~ @q ~O�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~�^sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�asq ~�vsq ~�{q ~ �sq ~�}q ~�dsq ~�vsq ~�{q ~ �sq ~�}q ~�gsq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�lsq ~��uq ~��   q ~�lsq ~��sq ~��?@     q ~�lq ~�gxq ~�guq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�gxq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~�vsq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�{sq ~��uq ~��   sq ~��uq ~��   q ~�{sq ~��sq ~��?@     q ~�aq ~�{xq ~�auq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�{q ~�vsq ~��sq ~��?@     q ~�vq ~�dq ~�{xq ~�duq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~�vq ~�aq ~�dq ~�{xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�aq ~�vq ~�dxq ~ �q ~��q ~	!uq ~��   q ~ �q ~sq ~��sq ~��?@     q ~�dq ~�axq ~Jsq ~��sq ~��?@     q ~�gq ~�aq ~�dxq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~�dq ~�axq ~	,sq ~��sq ~��?@     q ~�axq ~�q ~��q ~���sq ~��='S   sq ~���w��   sq ~���ƥ�   q ~�	q ~��q ~��sq ~���P�   q ~�q ~�	q ~��q ~��q ~��q ~��w   ;sq ~�gs�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~9sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~Euq ~��   q ~ �q ~Jq ~ <q ~��q ~	,�n��sq ~���ƥY   q ~�	q ~��q ~��w   sq ~�g����sq ~ sq ~ sq ~ 
w   q ~�<xq ~��q ~��sq ~ @q ~$�sq ~ G���    sq ~ sq ~ J   w   q ~�xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��xq ~$�uq ~��   q ~ <q ~ <q ~ �q ~��q ~�<uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~ � ��~sq ~���P�   q ~�q ~�	q ~��w   !sq ~�g���sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~�3���sq ~���g�   sq ~���z�z   q ~��q ~��q ~��q ~��q ~��w   2sq ~�g�E�"sq ~ sq ~ sq ~ 
w   q ~�<xq ~�q ~�sq ~ @q ~jsq ~ G���    sq ~ sq ~ J   w   q ~�xq ~�sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�	sq ~�vsq ~�{q ~ <sq ~�}q ~�sq ~��uq ~��   sq ~��uq ~��   q ~�sq ~��sq ~��?@     q ~�q ~�	xq ~�	uq ~��   q ~ <q ~ �q ~�q ~�<uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~�	xq ~ �q ~��q ~��!d��sq ~��mLߍ   sq ~��ȠU�   q ~��q ~�	q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��w   sq ~�gK��"sq ~ sq ~ sq ~ 
w   q ~�<xq ~�q ~�sq ~ @q ~�4sq ~ G���    sq ~ sq ~ J   w   q ~�xq ~�"sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�%sq ~�vsq ~�{q ~ <sq ~�}q ~�(sq ~��uq ~��   sq ~��uq ~��   q ~�(sq ~��sq ~��?@     q ~�(q ~�%xq ~�%uq ~��   q ~ <q ~ �q ~�.q ~�<uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~�%xq ~ �q ~��q ~�ʁ�sq ~���9�   q ~�q ~�q ~��w   Asq ~�g����sq ~ sq ~ sq ~ 
w   q ~��q ~�xq ~�8q ~�7sq ~ @q ~sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~�<sq ~�qsq ~�vq ~��sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~��uq ~��   q ~ �q ~q ~ <q ~��q ~	,Z`O�q ~��w   sq ~�g��)sq ~ sq ~ sq ~ 
w   q ~��q ~�7xq ~�Iq ~�Hsq ~ @q ~�sq ~ G���    sq ~ sq ~ J   w   q ~	,q ~ <xq ~�Msq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~�7q ~��q ~Auq ~��   q ~q ~q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~����@q ~��w   Osq ~�gG0�Hsq ~ sq ~ sq ~ 
w   q ~�xq ~�\q ~�[sq ~ @q ~$�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�`sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��xq ~�uq ~��   q ~ <q ~ <q ~ �q ~�hq ~�uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~ �Fx��q ~��w   Hsq ~�g�+9Tsq ~ sq ~ sq ~ 
w   q ~�xq ~�qq ~�psq ~ @q ~W�sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~�usq ~�qsq ~�vsq ~�{q ~sq ~�}q ~�xsq ~�vsq ~�{q ~ �sq ~�}q ~�{sq ~�vsq ~�{q ~ �sq ~�}q ~�~sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~�{q ~��xq ~�{uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~�~q ~��xq ~�~uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�~q ~�{q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�~q ~�{xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~Euq ~��   q ~ �q ~Jq ~ <sq ~��sq ~��?@     q ~�{xq ~	,q ~��q ~�sq ~��sq ~��?@      xq ~���&`(sq ~���]�   sq ~���ƥY   q ~�	q ~��q ~��q ~�q ~��w   Lsq ~�g�n9sq ~ sq ~ sq ~ 
w   q ~��q ~�xq ~��q ~��sq ~ @q ~nsq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~��sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��xq ~	,q ~��q ~�sq ~��sq ~��?@      xq ~�iw�Aq ~�w   >sq ~�g�L(�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~Lsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~�qsq ~�vq ~� sq ~�vq ~�#sq ~��uq ~��   q ~�>sq ~��uq ~��   q ~� q ~�!q ~Huq ~��   q ~ :q ~sq ~��sq ~��?@     q ~�#q ~� xq ~Auq ~��   q ~q ~q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ ��GOaq ~�2w   #sq ~�g,���sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~��,���sq ~���9�   q ~�q ~�q ~��w    sq ~�g�؏�sq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @q ~sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vq ~��sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ �q ~q ~��q ~Jq ~��q ~��uq ~��   q ~ �q ~q ~ <q ~��q ~	,TXq ~��w   sq ~�gT��!sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~� sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~1vq ~��q ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~��S�0�q ~��w   sq ~�g���sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @q ~ �sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�sq ~�qsq ~�vq ~�@sq ~�vq ~�Csq ~��uq ~��   sq ~��uq ~��   q ~�Cq ~ �q ~�Dq ~�uq ~��   q ~ <q ~ <q ~ �q ~�Jsq ~��sq ~��?@     q ~�Cq ~�@xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�@xq ~ �q ~��q ~���Iq ~�Tw   +sq ~�g�[Bsq ~ sq ~ sq ~ 
w   q ~�xq ~�$q ~�#sq ~ @q ~nsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~�(sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~�uq ~��   q ~ �q ~Jq ~ <sq ~��sq ~��?@     q ~��xq ~	,q ~��q ~�sq ~��sq ~��?@      xq ~�˨�q ~�w   Gsq ~�g���Ssq ~ sq ~ sq ~ 
w   q ~��xq ~�;q ~�:sq ~ @q ~-sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�?sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~�q ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~sq ~��sq ~��?@     q ~��q ~��q ~��xq ~Euq ~��   q ~ �q ~Jq ~ <sq ~��sq ~��?@     q ~��q ~��xq ~	,sq ~��sq ~��?@     q ~��xq ~�q ~��q ~��
�_q ~�w   9sq ~�g�P3�sq ~ sq ~ sq ~ 
w    xq ~�Vq ~�Usq ~ @q ~�Isq ~ G  �    sq ~ sq ~ J    w    xq ~�Zsq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�]sq ~�vsq ~�{q ~ �sq ~�}q ~�`sq ~�vsq ~�{q ~ <sq ~�}q ~�csq ~��uq ~��   sq ~��uq ~��   q ~�csq ~��sq ~��?@     q ~�]q ~�cxq ~�]uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�csq ~��sq ~��?@     q ~�`q ~�cxq ~�`uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�`q ~�]q ~�cxq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�]q ~�`xq ~ �sq ~��sq ~��?@     q ~�]xq ~��q ~��q ~�3�P/�sq ~��8���   sq ~���k�   q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��q ~��q ~��w   
sq ~�gI�Ssq ~ sq ~ sq ~ 
w   q ~��xq ~�~q ~�}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ <sq ~��sq ~��?@     q ~��xq ~sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��xq ~Vq ~��q ~T�a�sq ~������   sq ~���ƥY   q ~�	q ~��q ~��q ~��q ~��w   $sq ~�g��B�sq ~ sq ~ sq ~ 
w   q ~�q ~��q ~�7xq ~��q ~��sq ~ @q ~�sq ~ G)���    sq ~ sq ~ J   w   q ~ �q ~	,q ~ <xq ~��sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��q ~��uq ~��   q ~ �q ~ <q ~�7q ~��q ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~��B��q ~��w   Qsq ~�g4W��sq ~ sq ~ sq ~ 
w   q ~��q ~��xq ~��q ~��sq ~ @q ~�sq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��xq ~ �q ~��q ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~	,sq ~��sq ~��?@     q ~��xq ~�q ~��q ~�[�B�sq ~���<�   sq ~����;!   sq ~���ƥ�   q ~�	q ~��q ~��sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��q ~��q ~��q ~��w   8sq ~�gk�ƹsq ~ sq ~ sq ~ 
w   q ~��q ~�xq ~�q ~�sq ~ @q ~W�sq ~ G�C�j    sq ~ sq ~ J   w   q ~Tq ~xq ~�sq ~�qsq ~�vq ~�xsq ~�vq ~�{sq ~�vq ~�~sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~q ~��q ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~�{xq ~	,q ~��q ~�sq ~��sq ~��?@      xq ~��7!�q ~��w   Bsq ~�gq�*�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @q ~@�sq ~ G  �    sq ~ sq ~ J    w    xq ~�#sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�&sq ~�vsq ~�{q ~ <sq ~�}q ~�)sq ~��uq ~��   q ~�)sq ~��sq ~��?@     q ~�&q ~�)xq ~�&uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�&xq ~ �q ~��q ~��q�'sq ~��	f�   q ~�sq ~��ȠU�   q ~��q ~�	q ~��q ~��w   .sq ~�g�[sq ~ sq ~ sq ~ 
w   q ~�xq ~�7q ~�6sq ~ @q ~��sq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~�;sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~�>sq ~��uq ~��   q ~�>q ~�?q ~�uq ~��   q ~ <q ~ <q ~��q ~jVB�sq ~����!�   q ~�	q ~�	q ~��w   sq ~�gYY�Qsq ~ sq ~ sq ~ 
w   q ~��xq ~�Gq ~�Fsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�Msq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�Psq ~�vsq ~�{q ~ �sq ~�}q ~�Ssq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�Xsq ~��uq ~��   sq ~��uq ~��   q ~�Xsq ~��sq ~��?@     q ~�Pq ~�Xxq ~�Puq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�Xsq ~��sq ~��?@     q ~�Sq ~�Xxq ~�Suq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�Pq ~�Sq ~�Xxq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�Sq ~�Pxq ~ �q ~�iq ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~�Pxq ~	,q ~��q ~�n�]sq ~��8���   sq ~���k�   q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��q ~��q ~��w   sq ~�g(W~sq ~ sq ~ sq ~ 
w    xq ~�tq ~�ssq ~ @q ~0�sq ~ G  �    sq ~ sq ~ J    w    xq ~�xsq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�{sq ~�vsq ~�{q ~ <sq ~�}q ~�~sq ~��uq ~��   q ~�~sq ~��sq ~��?@     q ~�{q ~�~xq ~�{uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�{xq ~ �q ~��q ~��(S�sq ~���z�M   q ~��q ~��q ~��w   sq ~�g�h��sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��q ~��q ~��q ~�h�sq ~����!�   q ~�	q ~�	q ~��w   sq ~�gÏn�sq ~ sq ~ sq ~ 
w   q ~��q ~��xq ~��q ~��sq ~ @q ~u�sq ~ G���    sq ~ sq ~ J   w   q ~Tq ~	,xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~��q ~��xq ~ �q ~��q ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~sq ~��sq ~��?@     q ~��q ~��q ~��xq ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~	,sq ~��sq ~��?@     q ~��xq ~�q ~��q ~��.-�sq ~��='S   sq ~���w��   sq ~���ƥ�   q ~�	q ~��q ~��sq ~���P�   q ~�q ~�	q ~��q ~��q ~��q ~��w   Jsq ~�g��Ysq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @q ~W�sq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vq ~�xsq ~�vq ~�{sq ~�vq ~�~sq ~��uq ~��   q ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~��q ~5uq ~��   q ~ :q ~q ~��q ~Jq ~��q ~��uq ~��   q ~ �q ~q ~ <sq ~��sq ~��?@     q ~�{xq ~	,q ~��q ~�sq ~��sq ~��?@      xq ~���#R�q ~��w   "sq ~�gIJ�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t #0tt #0t:txq ~��q ~��sq ~ @q ~` sq ~ G  T    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~� q ~��sq ~��sq ~��?@      xq ~ �
��ksq ~��ȠU�   q ~��q ~�	q ~��w   Nsq ~�gq�%{sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�sq ~�vsq ~�{q ~ <sq ~�}q ~�sq ~��uq ~��   q ~�sq ~��sq ~��?@     q ~�q ~�xq ~�uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�xq ~ �q ~��q ~��q�!�sq ~��	aJ   q ~�sq ~��ȠU�   q ~��q ~�	q ~��q ~��w   sq ~�g8/[�sq ~ sq ~ sq ~ 
w   q ~��xq ~�"q ~�!sq ~ @q ~	'sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�&sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�)sq ~�vsq ~�{q ~ �sq ~�}q ~�,sq ~�vsq ~�{q ~ �sq ~�}q ~�/sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�4sq ~��uq ~��   q ~�4sq ~��sq ~��?@     q ~�4q ~�/xq ~�/uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�/xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~�>sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�Csq ~��uq ~��   sq ~��uq ~��   q ~�Csq ~��sq ~��?@     q ~�)q ~�Cxq ~�)uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�Cq ~�>sq ~��sq ~��?@     q ~�>q ~�,q ~�Cxq ~�,uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~�)q ~�>q ~�,q ~�Cxq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�)q ~�>q ~�,xq ~ �q ~�Tq ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~�)q ~�,xq ~sq ~��sq ~��?@     q ~�)q ~�/q ~�,xq ~�uq ~��   q ~ �q ~Jq ~ <sq ~��sq ~��?@     q ~�)q ~�,xq ~	,sq ~��sq ~��?@     q ~�)xq ~�q ~��q ~�M^�sq ~��='S   sq ~���w��   sq ~���ƥ�   q ~�	q ~��q ~��sq ~���P�   q ~�q ~�	q ~��q ~��q ~��q ~��w   :sq ~�g@�H�sq ~ sq ~ sq ~ 
w   q ~�7xq ~�gq ~�fsq ~ @q ~Qsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�ksq ~�q ~�79|vq ~�	w   Tsq ~�gL�Zsq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~�pq ~�osq ~ @q ~Lsq ~ G�W9J    sq ~ sq ~ J   w   q ~ �q ~xq ~�tsq ~�qsq ~�vq ~� sq ~�vq ~�#sq ~��uq ~��   sq ~��uq ~��   q ~�#q ~�$q ~Huq ~��   q ~ :q ~q ~�Asq ~��sq ~��?@     q ~�#q ~� xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ �Ċ��q ~�2w   Ssq ~�gʆ�sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~��q ~��sq ~ @q ~Lsq ~ G�W9J    sq ~ sq ~ J   w   q ~ �q ~xq ~��sq ~�qsq ~�vq ~� sq ~�vq ~�#sq ~��uq ~��   q ~�>q ~��sq ~��sq ~��?@     q ~�#q ~� xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ �mG��q ~�2w   Psq ~�g���sq ~ sq ~ sq ~ 
w   q ~�q ~�7xq ~��q ~��sq ~ @q ~ �sq ~ G��S    sq ~ sq ~ J   w   q ~ �q ~ <xq ~��sq ~�qsq ~�vq ~�@sq ~�vq ~�Csq ~��uq ~��   sq ~��uq ~��   q ~�Cq ~�7q ~�Dq ~�uq ~��   q ~ <q ~ <q ~ �q ~�Jsq ~��sq ~��?@     q ~�Cq ~�@xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�@xq ~ �q ~��q ~��Z�Iq ~�Tw   Isq ~�g~W�sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @q ~O�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~	,sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~��xq ~	,q ~��sq ~ ��~t <<<e,t>,e>,<<e,t>,e>>q ~	,q ~	,~W�!sq ~�����z   sq ~���ƥ�   q ~�	q ~��q ~��sq ~���ƥY   q ~�	q ~��q ~��q ~��w   sq ~�g�	�@sq ~ sq ~ sq ~ 
w   q ~�<q ~�xq ~��q ~��sq ~ @q ~$�sq ~ G�Uܘ    sq ~ sq ~ J   w   q ~�q ~ �xq ~��sq ~�qsq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   sq ~��uq ~��   q ~��q ~��sq ~��sq ~��?@     q ~��q ~��xq ~�uq ~��   q ~ <q ~ <q ~ �q ~��q ~�<uq ~��   q ~ �q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~ �_p�q ~��w   Rsq ~�g��p�sq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~�sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�	sq ~��uq ~��   sq ~��uq ~��   q ~�	sq ~��sq ~��?@     q ~�	q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�	q ~�sq ~��sq ~��?@     q ~��q ~�	q ~�xq ~��uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~��q ~�	q ~��q ~�xq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~��q ~�q ~��xq ~ �q ~�q ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~��q ~��xq ~sq ~��sq ~��?@     q ~��q ~��q ~��xq ~�uq ~��   q ~ �q ~Jq ~ <sq ~��sq ~��?@     q ~��q ~��xq ~	,sq ~��sq ~��?@     q ~��xq ~�q ~��q ~��&��sq ~���<�   sq ~����;!   sq ~���ƥ�   q ~�	q ~��q ~��sq ~��(Iɟ   sq ~��ȠU�   q ~��q ~�	q ~��q ~�	q ~��q ~��q ~��q ~��w   Esq ~�gs>3qsq ~ sq ~ sq ~ 
w   q ~��xq ~�.q ~�-sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�4sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�7sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�<sq ~��uq ~��   q ~�<sq ~��sq ~��?@     q ~�<q ~�7xq ~�7uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�7xq ~ �q ~�Cq ~��uq ~��   q ~ �q ~ <q ~��q ~	,�m�}sq ~���ƥY   q ~�	q ~��q ~��w   sq ~�g��v�sq ~ sq ~ sq ~ 
w    xq ~�Jq ~�Isq ~ @q ~s�sq ~ G  �    sq ~ sq ~ J    w    xq ~�Nsq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�Qsq ~�vsq ~�{q ~ <sq ~�}q ~�Tsq ~��uq ~��   q ~�Tsq ~��sq ~��?@     q ~�Qq ~�Txq ~�Quq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�Qxq ~ �q ~��q ~�ʇ�r�sq ~��(J�]   sq ~��ȠU�   q ~��q ~�	q ~��q ~�q ~��w   sq ~�g�^�sq ~ sq ~ sq ~ 
w   q ~�7xq ~�bq ~�asq ~ @q ~�sq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�fsq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~�7q ~��q ~Auq ~��   q ~q ~q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~�����|q ~��w   Ksq ~�g���sq ~ sq ~ sq ~ 
w   q ~��xq ~�uq ~�tsq ~ @q ~�sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�ysq ~�qsq ~�vq ~��sq ~�vq ~��sq ~�vq ~��sq ~��uq ~��   q ~��q ~1vq ~��q ~Auq ~��   q ~q ~q ~ �sq ~��sq ~��?@     q ~��q ~��xq ~ �sq ~��sq ~��?@     q ~��xq ~��q ~��q ~��	�i(q ~��w   Fsq ~�g�O�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~�uq ~��   q ~ <q ~ <q ~��q ~fv�sq ~��ȠU�   q ~��q ~�	q ~��w   5sq ~�g���sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @q ~�sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��q ~��q ~��q ~����sq ~���|�   q ~��q ~��q ~��w   /sq ~�g�ҀQsq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ GW�m�    sq ~ sq ~ J   w   q ~Txq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��sq ~��sq ~��?@     q ~��q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~5uq ~��   q ~ :q ~q ~��q ~Jq ~��q ~��uq ~��   q ~ �q ~q ~ <q ~��q ~	,dQ�sq ~���ƥY   q ~�	q ~��q ~��w   sq ~�g>�#sq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @q ~O�sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~��sq ~�qsq ~�vq ~�asq ~�vq ~�dsq ~�vq ~�gsq ~��uq ~��   q ~�ksq ~�vq ~�vsq ~��uq ~��   q ~�zq ~��q ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~�dq ~�axq ~sq ~��sq ~��?@     q ~�gq ~�aq ~�dxq ~Euq ~��   q ~ �q ~Jq ~ <sq ~��sq ~��?@     q ~�dq ~�axq ~	,sq ~��sq ~��?@     q ~�axq ~�q ~��q ~�SBl/q ~��w   sq ~�gjw�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~Lsq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�qsq ~�vq ~� sq ~�vq ~�#sq ~��uq ~��   q ~�zq ~��sq ~��sq ~��?@     q ~�#q ~� xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ ���q ~�2w   1sq ~�g���^sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @q ~{sq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~��sq ~�vsq ~�{q ~ <sq ~�}q ~� sq ~��uq ~��   q ~� sq ~��sq ~��?@     q ~� q ~��xq ~��uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~��xq ~ �q ~��q ~�����~sq ~��mL1-   sq ~��ȠU�   q ~��q ~�	q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��w   sq ~�g���sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ @q ~z�sq ~ G  �    sq ~ sq ~ J    w    xq ~�sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�q ~�q ~��q ~����sq ~���|��   q ~��q ~��q ~��w   %sq ~�gI�psq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @q ~,�sq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~� sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~�#sq ~�vsq ~�{q ~ <sq ~�}q ~�&sq ~��uq ~��   q ~�#q ~�&sq ~��sq ~��?@     q ~�#q ~�&xq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~�#xq ~ �q ~��q ~ �H�o�sq ~���P�   q ~�q ~�	q ~��w   	sq ~�gn�g@sq ~ sq ~ sq ~ 
w   q ~��xq ~�3q ~�2sq ~ @q ~��sq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�7sq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�:sq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�?sq ~��uq ~��   q ~�?sq ~��sq ~��?@     q ~�?q ~�:xq ~�:uq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�:xq ~ �q ~�Fq ~��uq ~��   q ~ �q ~ <q ~��q ~	,�#�Lsq ~���|�(   q ~��q ~��q ~��w   sq ~�gI�psq ~ sq ~ sq ~ 
w   q ~�xq ~�Mq ~�Lsq ~ @q ~Asq ~ G?z��    sq ~ sq ~ J   w   q ~ �xq ~�Qsq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~�Tsq ~�vsq ~�{q ~ <sq ~�}q ~�Wsq ~��uq ~��   q ~�Wq ~�Tsq ~��sq ~��?@     q ~�Wq ~�Txq ~�uq ~��   q ~ <q ~ <q ~ �sq ~��sq ~��?@     q ~�Txq ~ �q ~��q ~ �H�o�sq ~���P�   q ~�q ~�	q ~��w   sq ~�gYE�sq ~ sq ~ sq ~ 
w   q ~��xq ~�dq ~�csq ~ @q ~Vpsq ~ GI:�t    sq ~ sq ~ J   w   q ~	,xq ~�hsq ~�qsq ~�vsq ~�{q ~ �sq ~�}q ~�ksq ~�vsq ~�{q ~ �sq ~�}q ~�nsq ~��uq ~��   sq ~�vsq ~�{q ~ <sq ~�}q ~�ssq ~��uq ~��   sq ~��uq ~��   q ~�ssq ~��sq ~��?@     q ~�kq ~�sxq ~�kuq ~��   q ~ <q ~ �sq ~��uq ~��   q ~�ssq ~��sq ~��?@     q ~�nq ~�sxq ~�nuq ~��   q ~ <q ~ �sq ~��sq ~��?@     q ~�nq ~�kq ~�sxq ~��uq ~��   q ~ �q ~ �q ~ �sq ~��sq ~��?@     q ~�nq ~�kxq ~ �q ~��q ~��uq ~��   q ~ �q ~ <sq ~��sq ~��?@     q ~�kxq ~	,q ~��q ~�nu
�sq ~��8���   sq ~���f   q ~��sq ~��ȠU�   q ~��q ~�	q ~��q ~��q ~��q ~��w   (sq ~�g��sq ~ sq ~ sq ~ 
w    xq ~��q ~��sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~��sq ~�qsq ~�vsq ~�{q ~ <sq ~�}q ~��q ~��q ~��q ~���sq ~��ȠU�   q ~��q ~�	q ~��w   sq ~�g��'sq ~ sq ~ sq ~ 
w   q ~��xq ~��q ~��sq ~ @q ~n�sq ~ G|#    sq ~ sq ~ J   w   q ~ �xq ~��sq ~�sq ~�vsq ~�{q ~ <sq ~�}q ~��sq ~��uq ~��   q ~��q ~��q ~��uq ~��   q ~ <q ~ �q ~��q ~ ��Ǵq ~��w   sq ~�gG�sq ~ sq ~ sq ~ 
w   q ~�xq ~��q ~��sq ~ @q ~Lsq ~ G|!<    sq ~ sq ~ J   w   q ~xq ~��sq ~�qsq ~�vq ~� sq ~�vq ~�#sq ~��uq ~��   q ~�zq ~�Asq ~��sq ~��?@     q ~�#q ~� xq ~Auq ~��   q ~q ~q ~ �sq ~��sq ~��?@     q ~� xq ~ �q ~��q ~ ��h*q ~�2w   4xsq ~ !        sr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCoordinationFeatureSet�4tHWcg+ Z cpapFeaturesZ cpp1FeaturesZ reptFeaturesxpsr Dedu.cornell.cs.nlp.spf.parser.ccg.features.basic.RuleUsageFeatureSet�k�d�L2� D scaleZ unaryRulesOnlyL 	ignoreSetq ~ xp?������� sr java.util.HashSet�D�����4  xpw   ?@      xsr Ledu.cornell.cs.nlp.spf.parser.ccg.features.basic.DynamicWordSkippingFeatures%�q�� L emptyCategoryq ~�hL 
featureTagq ~ xpsq ~�p    sq ~��zT�lq ~��t EMPTYt DYNSKIPxq ~ sq ~ sq ~ J   w   q ~ xq ~��sr %java.util.Collections$UnmodifiableSet��я��U  xq ~ sq ~��w   ?@     sr .edu.cornell.cs.nlp.spf.base.hashvector.KeyArgs���]e.ɘ I hashCodeL arg1q ~ L arg2q ~ L arg3q ~ L arg4q ~ L arg5q ~ xp2Iݬq ~ t 
TMPDEFAULTpppsq ~��wzq ~ t XEMEDEFAULTpppsq ~��'��q ~ t 
LEXDEFAULTpppxsr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoredLexicon�>�"z L lexemesq ~ (L lexemesByTypeq ~ (L 	templatesq ~ (xpsq ~ C?@     w     -q ~L~sq ~��w   ?@     q ~Lsxq ~ sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�q ~�xq ~L�sq ~��w   ?@     q ~L�xq ~sq ~��w   ?@     q ~	xq ~�Bsq ~��w   ?@     q ~�7xq ~S2sq ~��w   ?@     q ~S'xq ~+ksq ~��w   ?@     q ~+`xq ~T�sq ~��w   ?@     q ~T�xq ~*hsq ~��w   ?@     q ~*]xq ~r�sq ~��w   ?@     q ~r�xq ~=�sq ~��w   ?@     q ~=�xq ~�sq ~��w   ?@     q ~�xq ~hVsq ~��w   ?@     q ~hKxq ~^sq ~��w   ?@     q ~Xxq ~��sq ~��w   ?@     q ~�vxq ~z�sq ~��w   ?@     q ~z�xq ~omsq ~��w   ?@     q ~o_q ~1�xq ~2%sq ~��w   ?@     q ~2q ~e�xq ~0�sq ~��w   ?@     q ~0�xq ~Zysq ~��w   ?@     q ~Znxq ~J�sq ~��w   ?@     q ~J�xq ~+�sq ~��w   ?@     q ~+�xq ~_Zsq ~��w   ?@     q ~_Oxq ~H�sq ~��w   ?@     q ~kvq ~H�xq ~3Qsq ~��w   ?@     q ~3Fxq ~#�sq ~��w   ?@     q ~#�xq ~DGsq ~��w   ?@     q ~[�q ~D<xq ~Vsq ~��w   ?@     q ~U�xq ~�sq ~��w   ?@     q ~cq ~�xq ~5sq ~��w   ?@     q ~5xq ~usq ~��w   ?@     q ~gq ~C�xq ~cTsq ~��w   ?@     q ~��q ~cIxq ~7�sq ~��w   ?@     q ~7txq ~1#sq ~��w   ?@     q ~1xq ~:�sq ~��w   ?@     q ~:�xq ~�sq ~��w   ?@     q ~�xq ~sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~`�sq ~��w   ?@     q ~pq ~`�xq ~��sq ~��w   ?@     q ~��q ~o|xq ~.Usq ~��w   ?@     q ~.Gxq ~)sq ~��w   ?@     q ~xq ~Ksq ~��w   ?@     q ~@xq ~J�sq ~��w   ?@     q ~J�xq ~�4sq ~��w   ?@     q ~�)xq ~�sq ~��w   ?@     q ~�xq ~%Jsq ~��w   ?@     q ~%?xq ~8sq ~��w   ?@     q ~8xq ~@jsq ~��w   ?@     q ~@_xq ~C$sq ~��w   ?@     q ~Cxq ~#sq ~��w   ?@     q ~"�q ~A�xq ~;sq ~��w   ?@     q ~0xq ~j�sq ~��w   ?@     q ~j�xq ~}�sq ~��w   ?@     q ~}�xq ~d:sq ~��w   ?@     q ~d/xq ~a�sq ~��w   ?@     q ~a�xq ~m"sq ~��w   ?@     q ~mq ~)exq ~g�sq ~��w   ?@     q ~g�xq ~/sq ~��w   ?@     q ~/xq ~W?sq ~��w   ?@     q ~W4xq ~�Ysq ~��w   ?@     q ~�Nxq ~B�sq ~��w   ?@     q ~Byxq ~Efsq ~��w   ?@     q ~E[q ~uQxq ~X9sq ~��w   ?@     q ~&�q ~X,xq ~$xsq ~��w   ?@     q ~$jxq ~gsq ~��w   ?@     q ~gxq ~k�sq ~��w   ?@     q ~Wmq ~k�xq ~vusq ~��w   ?@     q ~vjxq ~z�sq ~��w   ?@     q ~z�xq ~ZBsq ~��w   ?@     q ~Z7xq ~sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~Tsq ~��w   ?@     q ~Txq ~]�sq ~��w   ?@     q ~]�xq ~-�sq ~��w   ?@     q ~-�xq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~8sq ~��w   ?@     q ~8xq ~�sq ~��w   ?@     q ~Yq ~�xq ~R~sq ~��w   ?@     q ~Rsxq ~QUsq ~��w   ?@     q ~QJxq ~B�sq ~��w   ?@     q ~B�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�Sq ~�xq ~sq ~��w   ?@     q ~K�q ~xq ~c�sq ~��w   ?@     q ~c�xq ~E�sq ~��w   ?@     q ~Euxq ~-sq ~��w   ?@     q ~,�xq ~	sq ~��w   ?@     q ~	
xq ~Pwsq ~��w   ?@     q ~Plxq ~#sq ~��w   ?@     q ~NZq ~xq ~0�sq ~��w   ?@     q ~0�xq ~G,sq ~��w   ?@     q ~Gxq ~rsq ~��w   ?@     q ~dxq ~E�sq ~��w   ?@     q ~E�xq ~3Dsq ~��w   ?@     q ~39xq ~w�sq ~��w   ?@     q ~�q ~w�xq ~s�sq ~��w   ?@     q ~s�xq ~ Lsq ~��w   ?@     q ~ >xq ~_1sq ~��w   ?@     q ~_&xq ~90sq ~��w   ?@     q ~9%xq ~HJsq ~��w   ?@     q ~H?q ~3mxq ~�sq ~��w   ?@     q ~�q ~Q�xq ~X�sq ~��w   ?@     q ~X�q ~'�xq ~,$sq ~��w   ?@     q ~,xq ~~�sq ~��w   ?@     q ~~�xq ~��sq ~��w   ?@     q ~��q ~uxq ~t�sq ~��w   ?@     q ~t�xq ~(�sq ~��w   ?@     q ~(uxq ~(�sq ~��w   ?@     q ~(�xq ~hsq ~��w   ?@     q ~g�xq ~$sq ~��w   ?@     q ~$xq ~M�sq ~��w   ?@     q ~M�q ~d�xq ~�sq ~��w   ?@     q ~�xq ~)�sq ~��w   ?@     q ~)�xq ~�sq ~��w   ?@     q ~rxq ~.�sq ~��w   ?@     q ~.�xq ~Rsq ~��w   ?@     q ~Q�q ~Vxq ~B�sq ~��w   ?@     q ~B�xq ~	�sq ~��w   ?@     q ~	txq ~��sq ~��w   ?@     q ~�xq ~Rsq ~��w   ?@     q ~�sq ~Exq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�q ~q�xq ~��sq ~��w   ?@     q ~��xq ~A�sq ~��w   ?@     q ~A�q ~D-xq ~qssq ~��w   ?@     q ~qhxq ~$/sq ~��w   ?@     q ~$$xq ~��sq ~��w   ?@     q ~��xq ~crsq ~��w   ?@     q ~ceq ~�Uxq ~r�sq ~��w   ?@     q ~r�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~>�sq ~��w   ?@     q ~>�xq ~��sq ~��w   ?@     q ~��xq ~H�sq ~��w   ?@     q ~H�q ~�xq ~sq ~��w   ?@     q ~xq ~m�sq ~��w   ?@     q ~m�xq ~[8sq ~��w   ?@     q ~[+q ~G�xq ~0�sq ~��w   ?@     q ~0�xq ~Y)sq ~��w   ?@     q ~Yq ~�q ~IPxq ~.�sq ~��w   ?@     q ~.�xq ~��sq ~��w   ?@     q ~��q ~^/xq ~Sssq ~��w   ?@     q ~Shxq ~P]sq ~��w   ?@     q ~PRxq ~.(sq ~��w   ?@     q ~. xq ~z�sq ~��w   ?@     q ~z�xq ~}�sq ~��w   ?@     q ~}�xq ~)�sq ~��w   ?@     q ~)�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~vxq ~'(sq ~��w   ?@     q ~'xq ~[)sq ~��w   ?@     q ~[q ~zgxq ~ssq ~��w   ?@     q ~sxq ~3�sq ~��w   ?@     q ~3}xq ~�sq ~��w   ?@     q ~eq ~_�q ~xxq ~INsq ~��w   ?@     q ~ICxq ~ksq ~��w   ?@     q ~`q ~�xq ~(�sq ~��w   ?@     q ~(�xq ~lsq ~��w   ?@     q ~^xq ~I�sq ~��w   ?@     q ~I�xq ~��sq ~��w   ?@     q ~��xq ~>nsq ~��w   ?@     q ~>cxq ~��sq ~��w   ?@     q ~��xq ~+�sq ~��w   ?@     q ~+~xq ~�vsq ~��w   ?@     q ~�kxq ~O�sq ~��w   ?@     q ~��q ~,�q ~O�xq ~�bsq ~��w   ?@     q ~�Wxq ~^csq ~��w   ?@     q ~^Xxq ~�sq ~��w   ?@     q ~�xq ~d-sq ~��w   ?@     q ~d'xq ~79sq ~��w   ?@     q ~>�q ~7.xq ~C1sq ~��w   ?@     q ~C&xq ~!sq ~��w   ?@     q ~xq ~�sq ~��w   ?@     q ~�xq ~AIsq ~��w   ?@     q ~A;xq ~ �sq ~��w   ?@     q ~ �xq ~m�sq ~��w   ?@     q ~m�xq ~=�sq ~��w   ?@     q ~=�q ~�xq ~e�sq ~��w   ?@     q ~e�xq ~oCsq ~��w   ?@     q ~}�q ~j;q ~j}q ~�Hq ~raq ~0�q ~o8xq ~%Zsq ~��w   ?@     q ~%Lxq ~ sq ~��w   ?@     q ~sAq ~ xq ~4�sq ~��w   ?@     q ~4�xq ~+�sq ~��w   ?@     q ~!q ~+�xq ~�sq ~��w   ?@     q ~�yq ~��xq ~*�sq ~��w   ?@     q ~*�xq ~q$sq ~��w   ?@     q ~qxq ~y�sq ~��w   ?@     q ~y�xq ~;�sq ~��w   ?@     q ~;�xq ~/�sq ~��w   ?@     q ~/�xq ~%�sq ~��w   ?@     q ~%�xq ~f~sq ~��w   ?@     q ~fsxq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~osq ~��w   ?@     q ~n�q ~=}xq ~v>sq ~��w   ?@     q ~v0xq ~1osq ~��w   ?@     q ~1axq ~;�sq ~��w   ?@     q ~;�xq ~&�sq ~��w   ?@     q ~&�xq ~�1sq ~��w   ?@     q ~�&xq ~��sq ~��w   ?@     q ~�~xq ~�sq ~��w   ?@     q ~�xq ~Q�sq ~��w   ?@     q ~Q�xq ~!^sq ~��w   ?@     q ~!Sxq ~~sq ~��w   ?@     q ~~xq ~sq ~��w   ?@     q ~_�q ~�xq ~(ssq ~��w   ?@     q ~(hxq ~,�sq ~��w   ?@     q ~,�xq ~tsq ~��w   ?@     q ~ixq ~?sq ~��w   ?@     q ~>�xq ~��sq ~��w   ?@     q ~��xq ~�Psq ~��w   ?@     q ~�Exq ~E�sq ~��w   ?@     q ~E�xq ~pJsq ~��w   ?@     q ~p<q ~C3xq ~}�sq ~��w   ?@     q ~}�xq ~sq ~��w   ?@     q ~~Nq ~xq ~0sq ~��w   ?@     q ~"xq ~:Usq ~��w   ?@     q ~:Jxq ~R0sq ~��w   ?@     q ~Wq ~R#xq ~gsq ~��w   ?@     q ~\xq ~�sq ~��w   ?@     q ~�xq ~1�sq ~��w   ?@     q ~1�xq ~�sq ~��w   ?@     q ~�xq ~Osq ~��w   ?@     q ~N�xq ~Qsq ~��w   ?@     q ~P�xq ~4�sq ~��w   ?@     q ~4�xq ~�sq ~��w   ?@     q ~9�q ~�xq ~2nsq ~��w   ?@     q ~2cq ~,�xq ~��sq ~��w   ?@     q ~�vxq ~W]sq ~��w   ?@     q ~WNxq ~��sq ~��w   ?@     q ~��xq ~Rqsq ~��w   ?@     q ~Rfxq ~!1sq ~��w   ?@     q ~&�q ~!#xq ~|sq ~��w   ?@     q ~oxq ~�dsq ~��w   ?@     q ~�Yxq ~37sq ~��w   ?@     q ~3,xq ~0^sq ~��w   ?@     q ~0Pxq ~Y�sq ~��w   ?@     q ~Y�xq ~?�sq ~��w   ?@     q ~?�xq ~5Asq ~��w   ?@     q ~56xq ~g@sq ~��w   ?@     q ~g5xq ~�sq ~��w   ?@     q ~��xq ~@sq ~��w   ?@     q ~@	q ~xxq ~W�sq ~��w   ?@     q ~�q ~Wzxq ~�
sq ~��w   ?@     q ~��xq ~'Ysq ~��w   ?@     q ~'Kxq ~'�sq ~��w   ?@     q ~'�xq ~�sq ~��w   ?@     q ~��q ~C�xq ~bssq ~��w   ?@     q ~bexq ~o�sq ~��w   ?@     q ~o�xq ~TVsq ~��w   ?@     q ~TIxq ~}sq ~��w   ?@     q ~}xq ~6Xsq ~��w   ?@     q ~E�q ~6Jxq ~��sq ~��w   ?@     q ~�$q ~��xq ~usq ~��w   ?@     q ~jxq ~zesq ~��w   ?@     q ~zZxq ~�sq ~��w   ?@     q ~�xq ~k�sq ~��w   ?@     q ~k�xq ~j�sq ~��w   ?@     q ~#�q ~j�xq ~
-sq ~��w   ?@     q ~
xq ~(�sq ~��w   ?@     q ~(�q ~k(xq ~o�sq ~��w   ?@     q ~o�xq ~exsq ~��w   ?@     q ~emxq ~h�sq ~��w   ?@     q ~h�xq ~Z�sq ~��w   ?@     q ~Z�q ~T�xq ~:bsq ~��w   ?@     q ~:Wxq ~kgsq ~��w   ?@     q ~k\xq ~0�sq ~��w   ?@     q ~0�q ~Xxq ~�}sq ~��w   ?@     q ~�rxq ~Iksq ~��w   ?@     q ~I`xq ~�sq ~��w   ?@     q ~�q ~s�xq ~�sq ~��w   ?@     q ~yxq ~ltsq ~��w   ?@     q ~lfxq ~!�sq ~��w   ?@     q ~!�xq ~3sq ~��w   ?@     q ~3xq ~X�sq ~��w   ?@     q ~X�xq ~dsq ~��w   ?@     q ~c�xq ~[�sq ~��w   ?@     q ~[�xq ~"�sq ~��w   ?@     q ~"�xq ~4/sq ~��w   ?@     q ~4$xq ~0�sq ~��w   ?@     q ~0�xq ~(sq ~��w   ?@     q ~xq ~+
sq ~��w   ?@     q ~*�q ~=�xq ~l8sq ~��w   ?@     q ~l*xq ~f�sq ~��w   ?@     q ~f�xq ~Fsq ~��w   ?@     q ~Fxq ~x�sq ~��w   ?@     q ~x�q ~vxq ~�'sq ~��w   ?@     q ~�xq ~sq ~��w   ?@     q ~�xq ~S�sq ~��w   ?@     q ~S�xq ~9wsq ~��w   ?@     q ~9ixq ~�sq ~��w   ?@     q ~�xq ~q�sq ~��w   ?@     q ~q�xq ~H�sq ~��w   ?@     q ~H�q ~T�xq ~^�sq ~��w   ?@     q ~^�xq ~Mhsq ~��w   ?@     q ~MZxq ~�psq ~��w   ?@     q ~�exq ~N�sq ~��w   ?@     q ~N�xq ~,gsq ~��w   ?@     q ~,\xq ~Ysq ~��w   ?@     q ~qq ~�wq ~X�q ~Yq ~KRq ~M�xq ~=sq ~��w   ?@     q ~/q ~Y+xq ~T}sq ~��w   ?@     q ~Trxq ~ �sq ~��w   ?@     q ~ �q ~4�xq ~0 sq ~��w   ?@     q ~0xq ~h�sq ~��w   ?@     q ~hvq ~�xq ~gMsq ~��w   ?@     q ~gBxq ~(�sq ~��w   ?@     q ~(�xq ~3sq ~��w   ?@     q ~%xq ~�sq ~��w   ?@     q ~�xq ~|fsq ~��w   ?@     q ~|[xq ~7�sq ~��w   ?@     q ~7�xq ~�sq ~��w   ?@     q ~�q ~_dxq ~� sq ~��w   ?@     q ~��xq ~f�sq ~��w   ?@     q ~f�xq ~tesq ~��w   ?@     q ~i�q ~�>q ~@lq ~tZxq ~1sq ~��w   ?@     q ~1xq ~qLsq ~��w   ?@     q ~qAxq ~*:sq ~��w   ?@     q ~*/xq ~~ssq ~��w   ?@     q ~~hxq ~|Hsq ~��w   ?@     q ~|=xq ~qYsq ~��w   ?@     q ~qNxq ~�sq ~��w   ?@     q ~�xq ~v�sq ~��w   ?@     q ~v�xq ~�sq ~��w   ?@     q ~9�q ~�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�xq ~L#sq ~��w   ?@     q ~Lxq ~aRsq ~��w   ?@     q ~aGxq ~b<sq ~��w   ?@     q ~�q ~b/xq ~)�sq ~��w   ?@     q ~)�xq ~�sq ~��w   ?@     q ~�xq ~Yjsq ~��w   ?@     q ~Y_xq ~
sq ~��w   ?@     q ~
txq ~�sq ~��w   ?@     q ~�xq ~b sq ~��w   ?@     q ~�"q ~bq ~�Fxq ~9Wsq ~��w   ?@     q ~9Lq ~��xq ~\@sq ~��w   ?@     q ~\5q ~Yyxq ~Jsq ~��w   ?@     q ~<xq ~{$sq ~��w   ?@     q ~{xq ~K�sq ~��w   ?@     q ~K�xq ~f sq ~��w   ?@     q ~fxq ~��sq ~��w   ?@     q ~��xq ~sq ~��w   ?@     q ~xq ~y3sq ~��w   ?@     q ~y(xq ~�sq ~��w   ?@     q ~�xq ~a&sq ~��w   ?@     q ~axq ~ssq ~��w   ?@     q ~exq ~�sq ~��w   ?@     q ~�xq ~lsq ~��w   ?@     q ~lxq ~J`sq ~��w   ?@     q ~$q ~JSxq ~uBsq ~��w   ?@     q ~u7xq ~3�sq ~��w   ?@     q ~3�xq ~sq ~��w   ?@     q ~UJq ~xq ~�wsq ~��w   ?@     q ~�lxq ~#Fsq ~��w   ?@     q ~#;xq ~)�sq ~��w   ?@     q ~ _q ~)�xq ~sq ~��w   ?@     q ~xq ~(sq ~��w   ?@     q ~(xq ~oPsq ~��w   ?@     q ~oExq ~b�sq ~��w   ?@     q ~b�xq ~F�sq ~��w   ?@     q ~Fxq ~�sq ~��w   ?@     q ~��xq ~fdsq ~��w   ?@     q ~fYxq ~[�sq ~��w   ?@     q ~[�xq ~s�sq ~��w   ?@     q ~sxq ~d�q ~�xq ~%�sq ~��w   ?@     q ~%�xq ~f-sq ~��w   ?@     q ~f"xq ~�tsq ~��w   ?@     q ~�ixq ~��sq ~��w   ?@     q ~�~xq ~^�sq ~��w   ?@     q ~^�xq ~{�sq ~��w   ?@     q ~{~xq ~Psq ~��w   ?@     q ~O�xq ~s�sq ~��w   ?@     q ~'mq ~s�xq ~R�sq ~��w   ?@     q ~R�xq ~/�sq ~��w   ?@     q ~/txq ~�sq ~��w   ?@     q ~�xq ~)sq ~��w   ?@     q ~xq ~3�sq ~��w   ?@     q ~3�xq ~t�sq ~��w   ?@     q ~t�xq ~�sq ~��w   ?@     q ~^�q ~~xq ~+Nsq ~��w   ?@     q ~+@q ~1�xq ~Y�sq ~��w   ?@     q ~Y�xq ~sq ~��w   ?@     q ~�xq ~�-sq ~��w   ?@     q ~�"xq ~eZsq ~��w   ?@     q ~eOxq ~U�sq ~��w   ?@     q ~q ~U�xq ~/�sq ~��w   ?@     q ~/�xq ~�sq ~��w   ?@     q ~�xq ~'jsq ~��w   ?@     q ~'\xq ~E>sq ~��w   ?@     q ~E3xq ~h,sq ~��w   ?@     q ~h!xq ~��sq ~��w   ?@     q ~��xq ~5�sq ~��w   ?@     q ~5�xq ~sq ~��w   ?@     q ~xq ~/ sq ~��w   ?@     q ~/xq ~sq ~��w   ?@     q ~�xq ~;Tsq ~��w   ?@     q ~;Gq ~5�q ~Kixq ~]Ysq ~��w   ?@     q ~]Nxq ~S%sq ~��w   ?@     q ~Sxq ~��sq ~��w   ?@     q ~�{xq ~1sq ~��w   ?@     q ~#xq ~�sq ~��w   ?@     q ~�q ~Mxq ~-�sq ~��w   ?@     q ~-�xq ~AWsq ~��w   ?@     q ~ALxq ~y�sq ~��w   ?@     q ~y�xq ~d�sq ~��w   ?@     q ~d�xq ~�sq ~��w   ?@     q ~�xq ~Ksq ~��w   ?@     q ~=xq ~f�sq ~��w   ?@     q ~f�xq ~�sq ~��w   ?@     q ~zq ~xq ~!nsq ~��w   ?@     q ~!`xq ~W�sq ~��w   ?@     q ~W�xq ~�sq ~��w   ?@     q ~�q ~[�q ~mq ~�{q ~1rq ~=fq ~p�xq ~.psq ~��w   ?@     q ~.exq ~�sq ~��w   ?@     q ~�q ~�xq ~{Usq ~��w   ?@     q ~{Jxq ~z�sq ~��w   ?@     q ~^�q ~zwxq ~.�sq ~��w   ?@     q ~.�xq ~^Vsq ~��w   ?@     q ~^Kq ~ �xq ~;Dsq ~��w   ?@     q ~;6xq ~%�sq ~��w   ?@     q ~%�xq ~�rsq ~��w   ?@     q ~�q ~�gxq ~p�sq ~��w   ?@     q ~p�q ~*�xq ~�sq ~��w   ?@     q ~�xq ~k�sq ~��w   ?@     q ~k�xq ~��sq ~��w   ?@     q ~��q ~�@xq ~PCsq ~��w   ?@     q ~P8xq ~��sq ~��w   ?@     q ~��xq ~W�sq ~��w   ?@     q ~W�xq ~Vsq ~��w   ?@     q ~Hq ~K�xq ~a�sq ~��w   ?@     q ~a�xq ~~�sq ~��w   ?@     q ~~�xq ~��sq ~��w   ?@     q ~��xq ~H�sq ~��w   ?@     q ~2�q ~Hwxq ~'sq ~��w   ?@     q ~xq ~!�sq ~��w   ?@     q ~!�xq ~xusq ~��w   ?@     q ~xjxq ~ �sq ~��w   ?@     q ~ �xq ~�sq ~��w   ?@     q ~Z�q ~�xq ~��sq ~��w   ?@     q ~��xq ~*xsq ~��w   ?@     q ~*jxq ~ssq ~��w   ?@     q ~r�q ~tKxq ~%�sq ~��w   ?@     q ~%�q ~'�xq ~3�sq ~��w   ?@     q ~3�xq ~9�sq ~��w   ?@     q ~9�xq ~�fsq ~��w   ?@     q ~�[xq ~e�sq ~��w   ?@     q ~e�xq ~YPsq ~��w   ?@     q ~YExq ~*Isq ~��w   ?@     q ~*<xq ~l�sq ~��w   ?@     q ~l�xq ~Gsq ~��w   ?@     q ~Gxq ~sq ~��w   ?@     q ~�xq ~H�sq ~��w   ?@     q ~H�q ~0�xq ~C\sq ~��w   ?@     q ~CQxq ~S�sq ~��w   ?@     q ~S�xq ~'�sq ~��w   ?@     q ~a(q ~'�xq ~>�sq ~��w   ?@     q ~>yxq ~�=sq ~��w   ?@     q ~�2xq ~sq ~��w   ?@     q ~ xq ~�sq ~��w   ?@     q ~�q ~>xq ~P�sq ~��w   ?@     q ~Pyxq ~svsq ~��w   ?@     q ~skxq ~,�sq ~��w   ?@     q ~,�xq ~Ssq ~��w   ?@     q ~Exq ~u(sq ~��w   ?@     q ~uxq ~)�sq ~��w   ?@     q ~)rxq ~m�sq ~��w   ?@     q ~m�xq ~g�sq ~��w   ?@     q ~gvxq ~u�sq ~��w   ?@     q ~u�xq ~dksq ~��w   ?@     q ~d`q ~VNxq ~bVsq ~��w   ?@     q ~bKxq ~54sq ~��w   ?@     q ~5)xq ~ ]sq ~��w   ?@     q ~ Oxq ~Essq ~��w   ?@     q ~Ehxq ~T�sq ~��w   ?@     q ~T�xq ~�9sq ~��w   ?@     q ~�.xq ~��sq ~��w   ?@     q ~#�q ~��xq ~1�sq ~��w   ?@     q ~1�xq ~I�sq ~��w   ?@     q ~I�q ~�xq ~��sq ~��w   ?@     q ~��xq ~$�sq ~��w   ?@     q ~${xq ~3sq ~��w   ?@     q ~(xq ~3sq ~��w   ?@     q ~%xq ~[sq ~��w   ?@     q ~[xq ~�sq ~��w   ?@     q ~�q ~�#xq ~4�sq ~��w   ?@     q ~4�xq ~s?sq ~��w   ?@     q ~s4xq ~0�sq ~��w   ?@     q ~0�xq ~�
sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�xq ~|,sq ~��w   ?@     q ~|!xq ~�Xsq ~��w   ?@     q ~�Mxq ~��sq ~��w   ?@     q ~��xq ~"�sq ~��w   ?@     q ~"�xq ~H�sq ~��w   ?@     q ~H�xq ~�sq ~��w   ?@     q ~�xq ~Cvsq ~��w   ?@     q ~Ckxq ~��sq ~��w   ?@     q ~��xq ~�$sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��q ~<�xq ~h�sq ~��w   ?@     q ~#�q ~h�xq ~F�sq ~��w   ?@     q ~F�xq ~W�sq ~��w   ?@     q ~W�xq ~&rsq ~��w   ?@     q ~&dxq ~! sq ~��w   ?@     q ~ �xq ~:�sq ~��w   ?@     q ~:�xq ~|ssq ~��w   ?@     q ~|hxq ~�sq ~��w   ?@     q ~�xq ~ sq ~��w   ?@     q ~�xq ~xsq ~��w   ?@     q ~s�q ~xxq ~�sq ~��w   ?@     q ~|xq ~;nsq ~��w   ?@     q ~;cxq ~8�sq ~��w   ?@     q ~8�xq ~�.sq ~��w   ?@     q ~�#xq ~Asq ~��w   ?@     q ~@�xq ~"�sq ~��w   ?@     q ~"�xq ~G�sq ~��w   ?@     q ~Gzxq ~tsq ~��w   ?@     q ~txq ~x�sq ~��w   ?@     q ~x�q ~~!xq ~�
sq ~��w   ?@     q ~�xq ~u�sq ~��w   ?@     q ~u�xq ~�sq ~��w   ?@     q ~�xq ~htsq ~��w   ?@     q ~Eq ~hexq ~<Tsq ~��w   ?@     q ~<Gxq ~dzsq ~��w   ?@     q ~dmxq ~u�sq ~��w   ?@     q ~u�xq ~{Gsq ~��w   ?@     q ~{Aq ~~�xq ~jPsq ~��w   ?@     q ~jExq ~+sq ~��w   ?@     q ~xq ~I
sq ~��w   ?@     q ~H�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�q ~nxq ~�sq ~��w   ?@     q ~��q ~�xq ~|;sq ~��w   ?@     q ~~q ~|.xq ~>�sq ~��w   ?@     q ~>�xq ~S�sq ~��w   ?@     q ~S�xq ~�sq ~��w   ?@     q ~�xq ~W%sq ~��w   ?@     q ~Wxq ~+�sq ~��w   ?@     q ~+�q ~��xq ~U9sq ~��w   ?@     q ~U.xq ~�sq ~��w   ?@     q ~�xq ~hcsq ~��w   ?@     q ~hXxq ~(�sq ~��w   ?@     q ~(�xq ~Hdsq ~��w   ?@     q ~HYq ~1}xq ~g�sq ~��w   ?@     q ~wxq ~g�xq ~��sq ~��w   ?@     q ~��xq ~8�sq ~��w   ?@     q ~8�xq ~`sq ~��w   ?@     q ~`
xq ~Rdsq ~��w   ?@     q ~RYxq ~Ssq ~��w   ?@     q ~]q ~Exq ~u�sq ~��w   ?@     q ~u�xq ~Esq ~��w   ?@     q ~7xq ~b�sq ~��w   ?@     q ~b�xq ~N�sq ~��w   ?@     q ~N�q ~�qxq ~�/sq ~��w   ?@     q ~�$xq ~�sq ~��w   ?@     q ~Iq ~�xq ~��sq ~��w   ?@     q ~��q ~L�xq ~+�sq ~��w   ?@     q ~+�xq ~n�sq ~��w   ?@     q ~n�q ~b�xq ~R�sq ~��w   ?@     q ~R�xq ~*�sq ~��w   ?@     q ~*�xq ~�ysq ~��w   ?@     q ~�lq ~/xq ~ �sq ~��w   ?@     q ~ �xq ~;�sq ~��w   ?@     q ~;}xq ~-Gsq ~��w   ?@     q ~-9xq ~IAsq ~��w   ?@     q ~I6xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~'�sq ~��w   ?@     q ~'�xq ~
�sq ~��w   ?@     q ~
�xq ~'sq ~��w   ?@     q ~'xq ~S�sq ~��w   ?@     q ~S�q ~Hxq ~��sq ~��w   ?@     q ~[�q ~��xq ~"Fsq ~��w   ?@     q ~�q ~"8xq ~sq ~��w   ?@     q ~xq ~]ssq ~��w   ?@     q ~]hxq ~wsq ~��w   ?@     q ~qxq ~|�sq ~��w   ?@     q ~|�xq ~`tsq ~��w   ?@     q ~`ixq ~�sq ~��w   ?@     q ~�xq ~;$sq ~��w   ?@     q ~;xq ~;�sq ~��w   ?@     q ~;�xq ~;�sq ~��w   ?@     q ~;�xq ~��sq ~��w   ?@     q ~��q ~`�xq ~v�sq ~��w   ?@     q ~v�xq ~Qsq ~��w   ?@     q ~Qtxq ~ldsq ~��w   ?@     q ~lYxq ~Asq ~��w   ?@     q ~6xq ~I�sq ~��w   ?@     q ~I�xq ~(�sq ~��w   ?@     q ~(�xq ~n�sq ~��w   ?@     q ~xq ~n�q ~1�q ~c�xq ~*�sq ~��w   ?@     q ~*�xq ~/-sq ~��w   ?@     q ~/"q ~��xq ~W�sq ~��w   ?@     q ~W�xq ~Z�sq ~��w   ?@     q ~Z�xq ~1sq ~��w   ?@     q ~#xq ~/�sq ~��w   ?@     q ~/�xq ~M�sq ~��w   ?@     q ~M�xq ~=�sq ~��w   ?@     q ~=�xq ~wisq ~��w   ?@     q ~w^xq ~/Xsq ~��w   ?@     q ~/Mxq ~n>sq ~��w   ?@     q ~n3xq ~q�sq ~��w   ?@     q ~q�xq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�xq ~�csq ~��w   ?@     q ~�Xxq ~q�sq ~��w   ?@     q ~q�xq ~��sq ~��w   ?@     q ~��xq ~$�sq ~��w   ?@     q ~$�xq ~c�sq ~��w   ?@     q ~~�q ~c�xq ~VLsq ~��w   ?@     q ~�q ~V?xq ~s�sq ~��w   ?@     q ~s�xq ~fqsq ~��w   ?@     q ~ffxq ~B]sq ~��w   ?@     q ~BRxq ~��sq ~��w   ?@     q ~��xq ~q�sq ~��w   ?@     q ~q�xq ~�sq ~��w   ?@     q ~�xq ~V�sq ~��w   ?@     q ~}q ~V�xq ~��sq ~��w   ?@     q ~��q ~ixq ~h9sq ~��w   ?@     q ~h.xq ~8�sq ~��w   ?@     q ~8�xq ~�sq ~��w   ?@     q ~�xq ~z/sq ~��w   ?@     q ~z$xq ~�sq ~��w   ?@     q ~�xq ~a_sq ~��w   ?@     q ~aTxq ~8&sq ~��w   ?@     q ~8xq ~1�sq ~��w   ?@     q ~1�xq ~3 sq ~��w   ?@     q ~2�xq ~f�sq ~��w   ?@     q ~l:q ~f�xq ~cGsq ~��w   ?@     q ~c<xq ~K�sq ~��w   ?@     q ~K�xq ~y�sq ~��w   ?@     q ~yxxq ~?Bsq ~��w   ?@     q ~?7xq ~?�sq ~��w   ?@     q ~?�q ~6gxq ~Vsq ~��w   ?@     q ~Vxq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~Z�sq ~��w   ?@     q ~Z�xq ~��sq ~��w   ?@     q ~�yq ~�xq ~��sq ~��w   ?@     q ~��q ~Q�q ~p�xq ~H�sq ~��w   ?@     q ~H�xq ~��sq ~��w   ?@     q ~6tq ~��xq ~B�sq ~��w   ?@     q ~B�q ~5{q ~}�xq ~{
sq ~��w   ?@     q ~zKq ~z�xq ~JDsq ~��w   ?@     q ~J9xq ~�sq ~��w   ?@     q ~�xq ~esq ~��w   ?@     q ~exq ~�psq ~��w   ?@     q ~�cq ~�xq ~6�sq ~��w   ?@     q ~6�xq ~Xsq ~��w   ?@     q ~@q ~�q ~h�q ~x�xq ~9sq ~��w   ?@     q ~9xq ~K�sq ~��w   ?@     q ~K�xq ~c�sq ~��w   ?@     q ~c�xq ~�Zsq ~��w   ?@     q ~�Oxq ~��sq ~��w   ?@     q ~��xq ~qsq ~��w   ?@     q ~qxq ~<sq ~��w   ?@     q ~;�xq ~8�sq ~��w   ?@     q ~8wxq ~�sq ~��w   ?@     q ~�xq ~rsq ~��w   ?@     q ~rxq ~4rsq ~��w   ?@     q ~4gxq ~�lsq ~��w   ?@     q ~�_q ~Oxq ~Nsq ~��w   ?@     q ~@xq ~_�sq ~��w   ?@     q ~_�xq ~F�sq ~��w   ?@     q ~F�xq ~R�sq ~��w   ?@     q ~R�xq ~[sq ~��w   ?@     q ~[q ~��xq ~4!sq ~��w   ?@     q ~4xq ~_�sq ~��w   ?@     q ~_�q ~��xq ~_sq ~��w   ?@     q ~_xq ~�sq ~��w   ?@     q ~�xq ~
�sq ~��w   ?@     q ~
�q ~�xq ~}Gsq ~��w   ?@     q ~}<xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~>�sq ~��w   ?@     q ~rDq ~>�xq ~�jsq ~��w   ?@     q ~?�q ~�_xq ~5lsq ~��w   ?@     q ~5^xq ~B-sq ~��w   ?@     q ~B"q ~Mjxq ~-esq ~��w   ?@     q ~-Zxq ~`�sq ~��w   ?@     q ~`vq ~Q�xq ~d�sq ~��w   ?@     q ~d�xq ~%�sq ~��w   ?@     q ~%yxq ~>Esq ~��w   ?@     q ~>7xq ~Qsq ~��w   ?@     q ~Qxq ~B�sq ~��w   ?@     q ~B�xq ~SYsq ~��w   ?@     q ~SNxq ~��sq ~��w   ?@     q ~vMq ~��xq ~��sq ~��w   ?@     q ~��xq ~~�sq ~��w   ?@     q ~~�xq ~G
sq ~��w   ?@     q ~F�xq ~jsq ~��w   ?@     q ~i�xq ~\fsq ~��w   ?@     q ~\[xq ~�sq ~��w   ?@     q ~��xq ~(,sq ~��w   ?@     q ~(xq ~T*sq ~��w   ?@     q ~Txq ~=sq ~��w   ?@     q ~<�xq ~-rsq ~��w   ?@     q ~-gxq ~O�sq ~��w   ?@     q ~O�xq ~&Dsq ~��w   ?@     q ~&9q ~��xq ~�vsq ~��w   ?@     q ~�kxq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~g�sq ~��w   ?@     q ~;q ~g�xq ~5�sq ~��w   ?@     q ~5�xq ~\�sq ~��w   ?@     q ~\�xq ~Sfsq ~��w   ?@     q ~S[xq ~4�sq ~��w   ?@     q ~4�q ~{�xq ~g�sq ~��w   ?@     q ~g�xq ~-�sq ~��w   ?@     q ~-�xq ~�sq ~��w   ?@     q ~�xq ~g�sq ~��w   ?@     q ~g�xq ~�Dsq ~��w   ?@     q ~�9xq ~esq ~��w   ?@     q ~d�xq ~!�sq ~��w   ?@     q ~C�q ~!�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~;�q ~�xq ~m�sq ~��w   ?@     q ~m�xq ~l�sq ~��w   ?@     q ~l�q ~X xq ~�sq ~��w   ?@     q ~� xq ~N/sq ~��w   ?@     q ~N$xq ~`3sq ~��w   ?@     q ~`(xq ~v�sq ~��w   ?@     q ~v�xq ~ �sq ~��w   ?@     q ~ �xq ~,1sq ~��w   ?@     q ~,&xq ~8�sq ~��w   ?@     q ~q ~8�xq ~�7sq ~��w   ?@     q ~�,xq ~
Osq ~��w   ?@     q ~
Axq ~wvsq ~��w   ?@     q ~wkxq ~8�sq ~��w   ?@     q ~8�q ~M�xq ~C�sq ~��w   ?@     q ~C�xq ~*sq ~��w   ?@     q ~�q ~* xq ~?�sq ~��w   ?@     q ~?yxq ~j�sq ~��w   ?@     q ~j�xq ~kMsq ~��w   ?@     q ~kBxq ~>asq ~��w   ?@     q ~>Vxq ~�sq ~��w   ?@     q ~�xq ~[Usq ~��w   ?@     q ~[Gxq ~8usq ~��w   ?@     q ~8jxq ~}ysq ~��w   ?@     q ~}nxq ~E�sq ~��w   ?@     q ~E�xq ~$�sq ~��w   ?@     q ~$�q ~x[xq ~+�sq ~��w   ?@     q ~+�xq ~L�sq ~��w   ?@     q ~L�xq ~G�sq ~��w   ?@     q ~G�xq ~,�sq ~��w   ?@     q ~,vxq ~2Ssq ~��w   ?@     q ~2Exq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�xq ~,sq ~��w   ?@     q ~,xq ~o�sq ~��w   ?@     q ~o�xq ~1Rsq ~��w   ?@     q ~1Dxq ~hIsq ~��w   ?@     q ~h;xq ~GQsq ~��w   ?@     q ~GFxq ~V�sq ~��w   ?@     q ~V�xq ~&�sq ~��w   ?@     q ~&�xq ~osq ~��w   ?@     q ~axq ~6sq ~��w   ?@     q ~:q ~+xq ~fsq ~��w   ?@     q ~Yq ~B�xq ~'Hsq ~��w   ?@     q ~':xq ~:;sq ~��w   ?@     q ~:0xq ~x�sq ~��w   ?@     q ~�q ~x�xq ~}dsq ~��w   ?@     q ~}Yxq ~"sq ~��w   ?@     q ~!�xq ~�sq ~��w   ?@     q ~�xq ~<�sq ~��w   ?@     q ~<�xq ~~�sq ~��w   ?@     q ~~�xq ~�sq ~��w   ?@     q ~a�q ~�xq ~�Ksq ~��w   ?@     q ~�@xq ~]fsq ~��w   ?@     q ~][xq ~j9sq ~��w   ?@     q ~j.xq ~V�sq ~��w   ?@     q ~V�xq ~�0sq ~��w   ?@     q ~�"xq ~�>sq ~��w   ?@     q ~�3q ~U�xq ~6�sq ~��w   ?@     q ~6�q ~$�xq ~"sq ~��w   ?@     q ~xq ~'�sq ~��w   ?@     q ~'�xq ~H=sq ~��w   ?@     q ~H2xq ~�sq ~��w   ?@     q ~�xq ~N�sq ~��w   ?@     q ~N�xq ~dsq ~��w   ?@     q ~Vxq ~�sq ~��w   ?@     q ~�xq ~ktsq ~��w   ?@     q ~kixq ~P�sq ~��w   ?@     q ~P�xq ~=�sq ~��w   ?@     q ~=�q ~$]xq ~=�sq ~��w   ?@     q ~=�xq ~�sq ~��w   ?@     q ~�q ~oxq ~;sq ~��w   ?@     q ~-xq ~x-sq ~��w   ?@     q ~x"xq ~C�sq ~��w   ?@     q ~hq ~C�xq ~[sq ~��w   ?@     q ~Z�xq ~�sq ~��w   ?@     q ~�xq ~5�sq ~��w   ?@     q ~#q ~5�xq ~RWsq ~��w   ?@     q ~RLxq ~Tsq ~��w   ?@     q ~m�q ~S�xq ~#�sq ~��w   ?@     q ~#txq ~'�sq ~��w   ?@     q ~'�xq ~&�sq ~��w   ?@     q ~&�xq ~��sq ~��w   ?@     q ~Q�q ~��xq ~xsq ~��w   ?@     q ~mxq ~usq ~��w   ?@     q ~oq ~��xq ~W�sq ~��w   ?@     q ~W�xq ~�sq ~��w   ?@     q ~�xq ~� sq ~��w   ?@     q ~�xq ~3�sq ~��w   ?@     q ~3�xq ~0ksq ~��w   ?@     q ~0`q ~
�xq ~D�sq ~��w   ?@     q ~D�q ~2�xq ~>4sq ~��w   ?@     q ~>&xq ~5�sq ~��w   ?@     q ~5�xq ~/�sq ~��w   ?@     q ~/�xq ~]�sq ~��w   ?@     q ~]�xq ~d�sq ~��w   ?@     q ~d�xq ~|{sq ~��w   ?@     q ~|uxq ~"�sq ~��w   ?@     q ~"�xq ~"&sq ~��w   ?@     q ~"xq ~�sq ~��w   ?@     q ~rxq ~G�sq ~��w   ?@     q ~G�xq ~d$sq ~��w   ?@     q ~dxq ~"sq ~��w   ?@     q ~"
xq ~�qsq ~��w   ?@     q ~�fxq ~Ubsq ~��w   ?@     q ~UZxq ~)sq ~��w   ?@     q ~xq ~KCsq ~��w   ?@     q ~K8xq ~,sq ~��w   ?@     q ~xq ~�Zsq ~��w   ?@     q ~�Mq ~]'q ~�xq ~]�sq ~��w   ?@     q ~]uxq ~"�sq ~��w   ?@     q ~"�xq ~o6sq ~��w   ?@     q ~o+xq ~Ldsq ~��w   ?@     q ~LYxq ~9�sq ~��w   ?@     q ~9�xq ~ysq ~��w   ?@     q ~yq ~�xq ~+>sq ~��w   ?@     q ~+3xq ~P�sq ~��w   ?@     q ~P�xq ~�sq ~��w   ?@     q ~�q ~L�q ~xq ~N�sq ~��w   ?@     q ~Nvxq ~%sq ~��w   ?@     q ~xq ~^�sq ~��w   ?@     q ~^�xq ~F�sq ~��w   ?@     q ~F�xq ~%sq ~��w   ?@     q ~q ~x�xq ~:�sq ~��w   ?@     q ~:~xq ~BCsq ~��w   ?@     q ~B8xq ~�sq ~��w   ?@     q ~�xq ~\�sq ~��w   ?@     q ~\�xq ~F�sq ~��w   ?@     q ~F�xq ~�sq ~��w   ?@     q ~�q ~cxq ~nsq ~��w   ?@     q ~`xq ~m/sq ~��w   ?@     q ~m$xq ~Kgsq ~��w   ?@     q ~K\xq ~sq ~��w   ?@     q ~xq ~_�sq ~��w   ?@     q ~_�xq ~bcsq ~��w   ?@     q ~bXxq ~-�sq ~��w   ?@     q ~-�xq ~7rsq ~��w   ?@     q ~7jxq ~"�sq ~��w   ?@     q ~"�xq ~n�sq ~��w   ?@     q ~n�xq ~=Wsq ~��w   ?@     q ~=Iq ~yQxq ~Y�sq ~��w   ?@     q ~Y�xq ~��sq ~��w   ?@     q ~��xq ~M�sq ~��w   ?@     q ~Myxq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~��xq ~|�sq ~��w   ?@     q ~|~xq ~=sq ~��w   ?@     q ~=xq ~f�sq ~��w   ?@     q ~f�xq ~8gsq ~��w   ?@     q ~8Yxq ~x�sq ~��w   ?@     q ~x�xq ~1sq ~��w   ?@     q ~Doq ~+q ~Uxq ~,�sq ~��w   ?@     q ~,�xq ~esq ~��w   ?@     q ~Wq ~Fxq ~?jsq ~��w   ?@     q ~?\xq ~I{sq ~��w   ?@     q ~Imxq ~i�sq ~��w   ?@     q ~i}xq ~��sq ~��w   ?@     q ~7�q ~��xq ~J7sq ~��w   ?@     q ~J,q ~*xq ~{?sq ~��w   ?@     q ~{4xq ~�sq ~��w   ?@     q ~�q ~6�xq ~~�sq ~��w   ?@     q ~~�xq ~gZsq ~��w   ?@     q ~gOxq ~sq ~��w   ?@     q ~xq ~ dsq ~��w   ?@     q ~ Txq ~.csq ~��w   ?@     q ~.Xxq ~#9sq ~��w   ?@     q ~#+xq ~��sq ~��w   ?@     q ~aq ~��xq ~c�sq ~��w   ?@     q ~c�xq ~��sq ~��w   ?@     q ~��xq ~trsq ~��w   ?@     q ~tgxq ~|�sq ~��w   ?@     q ~|�xq ~ggsq ~��w   ?@     q ~g\xq ~h�sq ~��w   ?@     q ~h�q ~ lxq ~a�sq ~��w   ?@     q ~a�q ~N�xq ~Rsq ~��w   ?@     q ~0�q ~R
xq ~pdsq ~��w   ?@     q ~pYxq ~@�sq ~��w   ?@     q ~@{q ~T�xq ~0sq ~��w   ?@     q ~0xq ~y�sq ~��w   ?@     q ~y�xq ~d�sq ~��w   ?@     q ~q ~d�xq ~]sq ~��w   ?@     q ~Oxq ~�sq ~��w   ?@     q ~�xq ~gtsq ~��w   ?@     q ~gixq ~r_sq ~��w   ?@     q ~rTq ~E#xq ~6�sq ~��w   ?@     q ~6�xq ~#�sq ~��w   ?@     q ~#�xq ~"|sq ~��w   ?@     q ~"nxq ~D�sq ~��w   ?@     q ~D�xq ~��sq ~��w   ?@     q ~��xq ~Q�sq ~��w   ?@     q ~Q�xq ~6�sq ~��w   ?@     q ~6�xq ~��sq ~��w   ?@     q ~��xq ~M�sq ~��w   ?@     q ~M�xq ~1�sq ~��w   ?@     q ~pfq ~1�xq ~xsq ~��w   ?@     q ~ q ~mxq ~�sq ~��w   ?@     q ~�q ~�?xq ~a�sq ~��w   ?@     q ~a�xq ~]sq ~��w   ?@     q ~�q ~Oxq ~yvsq ~��w   ?@     q ~ykq ~Urxq ~&*sq ~��w   ?@     q ~&xq ~sq ~��w   ?@     q ~xq ~~�sq ~��w   ?@     q ~~�xq ~� sq ~��w   ?@     q ~�xq ~.�sq ~��w   ?@     q ~.�xq ~1sq ~��w   ?@     q ~1 xq ~Tpsq ~��w   ?@     q ~Texq ~GDsq ~��w   ?@     q ~G<xq ~,�sq ~��w   ?@     q ~w�q ~,�xq ~u�sq ~��w   ?@     q ~u{xq ~sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~?sq ~��w   ?@     q ~?q ~O#xq ~7	sq ~��w   ?@     q ~6�xq ~�sq ~��w   ?@     q ~�xq ~p�sq ~��w   ?@     q ~p�xq ~��sq ~��w   ?@     q ~��q ~Fxq ~h�sq ~��w   ?@     q ~h�xq ~	_sq ~��w   ?@     q ~	Qxq ~T:sq ~��w   ?@     q ~T,xq ~,sq ~��w   ?@     q ~+�xq ~�sq ~��w   ?@     q ~6�q ~�xq ~}sq ~��w   ?@     q ~|�xq ~11sq ~��w   ?@     q ~1&xq ~J*sq ~��w   ?@     q ~Jxq ~�jsq ~��w   ?@     q ~Qgq ~�\xq ~��sq ~��w   ?@     q ~��xq ~A�sq ~��w   ?@     q ~A�xq ~	�sq ~��w   ?@     q ~*�q ~	�xq ~Q�sq ~��w   ?@     q ~Q�xq ~�sq ~��w   ?@     q ~�xq ~Qsq ~��w   ?@     q ~t)q ~M�q ~<q ~eq ~F�xq ~8�sq ~��w   ?@     q ~8�xq ~*sq ~��w   ?@     q ~xq ~rsq ~��w   ?@     q ~rrq ~|�xq ~#�sq ~��w   ?@     q ~p�q ~#�xq ~r�sq ~��w   ?@     q ~r�xq ~	�sq ~��w   ?@     q ~	�xq ~&�sq ~��w   ?@     q ~&�xq ~�isq ~��w   ?@     q ~�^xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~J�sq ~��w   ?@     q ~J�q ~cVxq ~?Osq ~��w   ?@     q ~?Dxq ~#sq ~��w   ?@     q ~#q ~T�xq ~F�sq ~��w   ?@     q ~F�xq ~�sq ~��w   ?@     q ~�xq ~�Qsq ~��w   ?@     q ~�Fxq ~.�sq ~��w   ?@     q ~.�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~��q ~�xq ~�5sq ~��w   ?@     q ~�*xq ~Usq ~��w   ?@     q ~Jxq ~Wksq ~��w   ?@     q ~W`q ~l�xq ~c�sq ~��w   ?@     q ~w�q ~ctxq ~TGsq ~��w   ?@     q ~T<xq ~?(sq ~��w   ?@     q ~?xq ~$[sq ~��w   ?@     q ~$Pxq ~) sq ~��w   ?@     q ~(�xq ~I�sq ~��w   ?@     q ~I�xq ~uOsq ~��w   ?@     q ~uDxq ~[�sq ~��w   ?@     q ~[�xq ~A9sq ~��w   ?@     q ~A.xq ~n�sq ~��w   ?@     q ~n�xq ~{osq ~��w   ?@     q ~{dxq ~�7sq ~��w   ?@     q ~�,xq ~L�sq ~��w   ?@     q ~L�q ~B�xq ~�sq ~��w   ?@     q ~�xq ~p sq ~��w   ?@     q ~o�xq ~��sq ~��w   ?@     q ~��xq ~o�sq ~��w   ?@     q ~o�xq ~?sq ~��w   ?@     q ~1xq ~�sq ~��w   ?@     q ~[:q ~�xq ~,�sq ~��w   ?@     q ~,�xq ~O�sq ~��w   ?@     q ~O�q ~#�xq ~�sq ~��w   ?@     q ~�xq ~>Tsq ~��w   ?@     q ~>Gq ~axq ~)�sq ~��w   ?@     q ~)�xq ~M�sq ~��w   ?@     q ~M�xq ~7,sq ~��w   ?@     q ~7!xq ~h�sq ~��w   ?@     q ~h�xq ~R�sq ~��w   ?@     q ~R�q ~axq ~�sq ~��w   ?@     q ~�xq ~0Nsq ~��w   ?@     q ~t�q ~0@xq ~Ssq ~��w   ?@     q ~Exq ~X�sq ~��w   ?@     q ~X�xq ~S?sq ~��w   ?@     q ~S4xq ~9sq ~��w   ?@     q ~+xq ~	>sq ~��w   ?@     q ~	1q ~��xq ~sq ~��w   ?@     q ~)Xq ~	xq ~'�sq ~��w   ?@     q ~'~xq ~`�sq ~��w   ?@     q ~`�xq ~5�sq ~��w   ?@     q ~5�xq ~ysq ~��w   ?@     q ~kq ~}�xq ~^
sq ~��w   ?@     q ~]�xq ~X*sq ~��w   ?@     q ~Xxq ~��sq ~��w   ?@     q ~��xq ~_sq ~��w   ?@     q ~_xq ~8Vsq ~��w   ?@     q ~8Hxq ~�sq ~��w   ?@     q ~�xq ~Jsq ~��w   ?@     q ~]�q ~Jxq ~fsq ~��w   ?@     q ~fq ~a�xq ~/sq ~��w   ?@     q ~!xq ~`@sq ~��w   ?@     q ~`5xq ~Usq ~��w   ?@     q ~Jxq ~6;sq ~��w   ?@     q ~Gq ~6.xq ~�sq ~��w   ?@     q ~�xq ~G�sq ~��w   ?@     q ~G�xq ~7�sq ~��w   ?@     q ~7�xq ~9#sq ~��w   ?@     q ~9xq ~�5sq ~��w   ?@     q ~�*xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~zsq ~��w   ?@     q ~y�xq ~�sq ~��w   ?@     q ~�xq ~J�sq ~��w   ?@     q ~J�xq ~�csq ~��w   ?@     q ~�Xxq ~A+sq ~��w   ?@     q ~Axq ~^qsq ~��w   ?@     q ~^fxq ~�sq ~��w   ?@     q ~8(q ~�xq ~F}sq ~��w   ?@     q ~Frq ~�q ~xq ~sq ~��w   ?@     q ~�xq ~%�sq ~��w   ?@     q ~%�xq ~G:sq ~��w   ?@     q ~G/xq ~f�sq ~��w   ?@     q ~f�xq ~)=sq ~��w   ?@     q ~)/xq ~�sq ~��w   ?@     q ~�xq ~^-sq ~��w   ?@     q ~^"xq ~�Bsq ~��w   ?@     q ~�7xq ~�sq ~��w   ?@     q ~�xq ~R=sq ~��w   ?@     q ~R2xq ~D�sq ~��w   ?@     q ~D�q ~c�xq ~|�sq ~��w   ?@     q ~|�xq ~<�sq ~��w   ?@     q ~<�xq ~sq ~��w   ?@     q ~�xq ~\�sq ~��w   ?@     q ~\�xq ~[�sq ~��w   ?@     q ~[xq ~M�sq ~��w   ?@     q ~M�xq ~4sq ~��w   ?@     q ~3�q ~�xq ~b�sq ~��w   ?@     q ~b�xq ~]�sq ~��w   ?@     q ~]�xq ~2Csq ~��w   ?@     q ~28xq ~\�sq ~��w   ?@     q ~\uxq ~ksq ~��w   ?@     q ~aq ~kxq ~B�sq ~��w   ?@     q ~��q ~B�xq ~�Asq ~��w   ?@     q ~�6xq ~t�sq ~��w   ?@     q ~��q ~t�xq ~Usq ~��w   ?@     q ~Uxq ~,>sq ~��w   ?@     q ~,3xq ~&sq ~��w   ?@     q ~%�xq ~Fasq ~��w   ?@     q ~FVq ~oxq ~V�sq ~��w   ?@     q ~V�xq ~�sq ~��w   ?@     q ~�xq ~S�sq ~��w   ?@     q ~S}xq ~�sq ~��w   ?@     q ~�xq ~csq ~��w   ?@     q ~`Bq ~Vq ~dSxq ~�sq ~��w   ?@     q ~�q ~Y8xq ~~2sq ~��w   ?@     q ~~'xq ~P)sq ~��w   ?@     q ~Pxq ~i�sq ~��w   ?@     q ~i�xq ~msq ~��w   ?@     q ~mxq ~e sq ~��w   ?@     q ~exq ~Msq ~��w   ?@     q ~Mxq ~��sq ~��w   ?@     q ~��xq ~3*sq ~��w   ?@     q ~3q ~A�xq ~<sq ~��w   ?@     q ~1xq ~tIsq ~��w   ?@     q ~t>q ~�xq ~:�sq ~��w   ?@     q ~:�xq ~ �sq ~��w   ?@     q ~q ~tq ~\�q ~y5q ~ �xq ~isq ~��w   ?@     q ~ixq ~
�sq ~��w   ?@     q ~
�xq ~9sq ~��w   ?@     q ~9 xq ~�sq ~��w   ?@     q ~�q ~�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~xq ~�\sq ~��w   ?@     q ~�Qxq ~+^sq ~��w   ?@     q ~+Pq ~g�xq ~�sq ~��w   ?@     q ~�xq ~]�sq ~��w   ?@     q ~]�q ~y�xq ~sq ~��w   ?@     q ~_\q ~i>q ~xq ~1_sq ~��w   ?@     q ~1Txq ~ xsq ~��w   ?@     q ~ hxq ~=+sq ~��w   ?@     q ~= q ~x�xq ~
�sq ~��w   ?@     q ~
�q ~9Yxq ~m�sq ~��w   ?@     q ~m�xq ~hsq ~��w   ?@     q ~Zxq ~��sq ~��w   ?@     q ~�xxq ~T�sq ~��w   ?@     q ~T�xq ~V�sq ~��w   ?@     q ~V�xq ~k&sq ~��w   ?@     q ~kxq ~�sq ~��w   ?@     q ~�xq ~U�sq ~��w   ?@     q ~U�xq ~�sq ~��w   ?@     q ~�xq ~w�sq ~��w   ?@     q ~��q ~w�xq ~o�sq ~��w   ?@     q ~o�xq ~&asq ~��w   ?@     q ~&Sxq ~sq ~��w   ?@     q ~xq ~�esq ~��w   ?@     q ~�Zxq ~nsq ~��w   ?@     q ~v�q ~S�q ~nxq ~c:sq ~��w   ?@     q ~c/q ~�xq ~	.sq ~��w   ?@     q ~	q ~]�q ~p�xq ~Usq ~��w   ?@     q ~X;q ~��q ~Mxq ~Usq ~��w   ?@     q ~Gxq ~s�sq ~��w   ?@     q ~s�xq ~^�sq ~��w   ?@     q ~^�xq ~F�sq ~��w   ?@     q ~F�xq ~��sq ~��w   ?@     q ~��xq ~!�sq ~��w   ?@     q ~!�xq ~!�sq ~��w   ?@     q ~!�xq ~�sq ~��w   ?@     q ~zxq ~M6sq ~��w   ?@     q ~M(q ~Pxq ~:�sq ~��w   ?@     q ~:�q ~v�xq ~Bsq ~��w   ?@     q ~4xq ~r�sq ~��w   ?@     q ~r�xq ~:�sq ~��w   ?@     q ~:�xq ~Tcsq ~��w   ?@     q ~Mq ~TXxq ~O=sq ~��w   ?@     q ~O2xq ~|sq ~��w   ?@     q ~qxq ~O�sq ~��w   ?@     q ~N�q ~O�xq ~1Asq ~��w   ?@     q ~13xq ~}�sq ~��w   ?@     q ~}{xq ~/esq ~��w   ?@     q ~/Zq ~a8q ~v�xq ~=�sq ~��w   ?@     q ~=�xq ~/�sq ~��w   ?@     q ~/�xq ~��sq ~��w   ?@     q ~��q ~yDxq ~qfsq ~��w   ?@     q ~q[xq ~`�sq ~��w   ?@     q ~`�xq ~Y�sq ~��w   ?@     q ~Y�xq ~n�sq ~��w   ?@     q ~n�xq ~c�sq ~��w   ?@     q ~c�xq ~*-sq ~��w   ?@     q ~*q ~�xq ~%sq ~��w   ?@     q ~$�q ~P�q ~�"xq ~NKsq ~��w   ?@     q ~N>q ~Ixq ~��sq ~��w   ?@     q ~��q ~sxq ~_�sq ~��w   ?@     q ~_~xq ~�sq ~��w   ?@     q ~�xq ~C�sq ~��w   ?@     q ~C�xq ~��sq ~��w   ?@     q ~��xq ~`�sq ~��w   ?@     q ~`�xq ~4esq ~��w   ?@     q ~4Zq ~vwxq ~mVsq ~��w   ?@     q ~mKxq ~J�sq ~��w   ?@     q ~J�q ~Q0xq ~^�sq ~��w   ?@     q ~^�xq ~�Fsq ~��w   ?@     q ~�;xq ~	sq ~��w   ?@     q ~�xq ~n�sq ~��w   ?@     q ~n�xq ~ �sq ~��w   ?@     q ~ �xq ~o�sq ~��w   ?@     q ~o�xq ~'8sq ~��w   ?@     q ~'*xq ~]�sq ~��w   ?@     q ~]�xq ~Htsq ~��w   ?@     q ~Hnxq ~:sq ~��w   ?@     q ~,xq ~:sq ~��w   ?@     q ~:xq ~]�sq ~��w   ?@     q ~]�xq ~B sq ~��w   ?@     q ~Bxq ~�!sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~>�sq ~��w   ?@     q ~>�xq ~�sq ~��w   ?@     q ~�q ~xq ~z�sq ~��w   ?@     q ~z�xq ~R�sq ~��w   ?@     q ~R�q ~7xq ~v�sq ~��w   ?@     q ~v�xq ~
�sq ~��w   ?@     q ~
�xq ~fsq ~��w   ?@     q ~Xxq ~�sq ~��w   ?@     q ~�xq ~Zsq ~��w   ?@     q ~Zq ~g�xq ~esq ~��w   ?@     q ~Uxq ~N"sq ~��w   ?@     q ~Nq ~�xq ~sisq ~��w   ?@     q ~s^xq ~
sq ~��w   ?@     q ~
xq ~{bsq ~��w   ?@     q ~{Wxq ~X�sq ~��w   ?@     q ~X�xq ~3ksq ~��w   ?@     q ~3`xq ~d�sq ~��w   ?@     q ~�q ~d�xq ~7�sq ~��w   ?@     q ~7�xq ~:sq ~��w   ?@     q ~9�xq ~
�sq ~��w   ?@     q ~
�xq ~z<sq ~��w   ?@     q ~z1xq ~�sq ~��w   ?@     q ~�xq ~Ksq ~��w   ?@     q ~Kxq ~9�sq ~��w   ?@     q ~9�xq ~U�sq ~��w   ?@     q ~U�xq ~�sq ~��w   ?@     q ~9zq ~�xq ~�Usq ~��w   ?@     q ~�Oxq ~*Ysq ~��w   ?@     q ~*Kxq ~�sq ~��w   ?@     q ~�xq ~MFsq ~��w   ?@     q ~M8xq ~^�sq ~��w   ?@     q ~2q ~^�xq ~+{sq ~��w   ?@     q ~+mxq ~_Msq ~��w   ?@     q ~��q ~_@xq ~.sq ~��w   ?@     q ~.q ~�xq ~h�sq ~��w   ?@     q ~h�xq ~ �sq ~��w   ?@     q ~ yxq ~z�sq ~��w   ?@     q ~z�xq ~NXsq ~��w   ?@     q ~NMxq ~[�sq ~��w   ?@     q ~[�xq ~"lsq ~��w   ?@     q ~2q ~"axq ~��sq ~��w   ?@     q ~��xq ~usq ~��w   ?@     q ~gq ~H�xq ~v.sq ~��w   ?@     q ~v q ~�Rxq ~Nsq ~��w   ?@     q ~M�xq ~`Zsq ~��w   ?@     q ~`Oxq ~y�sq ~��w   ?@     q ~y�q ~�xq ~sq ~��w   ?@     q ~<Vq ~xq ~j�sq ~��w   ?@     q ~j�q ~	�xq ~M&sq ~��w   ?@     q ~Mxq ~@�sq ~��w   ?@     q ~@�xq ~a�sq ~��w   ?@     q ~Dyq ~a�xq ~Q�sq ~��w   ?@     q ~n_q ~Q�q ~6�xq ~EWsq ~��w   ?@     q ~EIxq ~$sq ~��w   ?@     q ~xq ~+�sq ~��w   ?@     q ~Hq ~+�xq ~[�sq ~��w   ?@     q ~[�xq ~^ sq ~��w   ?@     q ~[�q ~^xq ~u sq ~��w   ?@     q ~t�xq ~�sq ~��w   ?@     q ~�xq ~	Nsq ~��w   ?@     q ~	@q ~ZDxq ~"sq ~��w   ?@     q ~xq ~�<sq ~��w   ?@     q ~�1xq ~~Lsq ~��w   ?@     q ~~Axq ~l�sq ~��w   ?@     q ~l�xq ~w\sq ~��w   ?@     q ~wQxq ~X�sq ~��w   ?@     q ~X�xq ~�sq ~��w   ?@     q ~�xq ~5sq ~��w   ?@     q ~*xq ~hsq ~��w   ?@     q ~hxq ~!�sq ~��w   ?@     q ~!�xq ~&�sq ~��w   ?@     q ~[Xq ~&txq ~i"sq ~��w   ?@     q ~ixq ~O�sq ~��w   ?@     q ~O�xq ~0xsq ~��w   ?@     q ~0mxq ~K�sq ~��w   ?@     q ~K�xq ~�sq ~��w   ?@     q ~}fq ~�q ~u�xq ~Tsq ~��w   ?@     q ~Txq ~�sq ~��w   ?@     q ~-tq ~�xq ~W�sq ~��w   ?@     q ~W�xq ~K�sq ~��w   ?@     q ~�q ~K�xq ~�osq ~��w   ?@     q ~�dxq ~ Nsq ~��w   ?@     q ~ +xq ~usq ~��w   ?@     q ~uxq ~��sq ~��w   ?@     q ~��xq ~t<sq ~��w   ?@     q ~t1xq ~\&sq ~��w   ?@     q ~\xq ~ejsq ~��w   ?@     q ~e\xq ~gsq ~��w   ?@     q ~Zxq ~R�sq ~��w   ?@     q ~R�xq ~`�sq ~��w   ?@     q ~`�xq ~<"sq ~��w   ?@     q ~<xq ~G�sq ~��w   ?@     q ~G�xq ~dsq ~��w   ?@     q ~dq ~_xq ~Z*sq ~��w   ?@     q ~Zq ~x<xq ~|sq ~��w   ?@     q ~qxq ~b�sq ~��w   ?@     q ~b�xq ~#�sq ~��w   ?@     q ~#�xq ~��sq ~��w   ?@     q ~4q ~��xq ~x�sq ~��w   ?@     q ~x�xq ~G�sq ~��w   ?@     q ~G�q ~w�xq ~4�sq ~��w   ?@     q ~4�xq ~/Jsq ~��w   ?@     q ~/?xq ~r5sq ~��w   ?@     q ~*�q ~r(xq ~R�sq ~��w   ?@     q ~R�xq ~Usq ~��w   ?@     q ~Gxq ~��sq ~��w   ?@     q ~��xq ~Xsq ~��w   ?@     q ~Xyxq ~��sq ~��w   ?@     q ~��q ~p�xq ~�sq ~��w   ?@     q ~xxq ~�sq ~��w   ?@     q ~�xq ~$Msq ~��w   ?@     q ~aq ~$Bxq ~� sq ~��w   ?@     q ~�xq ~</sq ~��w   ?@     q ~<$xq ~?�sq ~��w   ?@     q ~?�xq ~��sq ~��w   ?@     q ~��xq ~z�sq ~��w   ?@     q ~z�xq ~V/sq ~��w   ?@     q ~V"q ~q'xq ~�sq ~��w   ?@     q ~�q ~Ngxq ~�sq ~��w   ?@     q ~�q ~
Sq ~xq ~r�sq ~��w   ?@     q ~r�xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~?�sq ~��w   ?@     q ~?�xq ~W�sq ~��w   ?@     q ~W�q ~7q ~�*q ~0xq ~J�sq ~��w   ?@     q ~Jxxq ~��sq ~��w   ?@     q ~��xq ~kZsq ~��w   ?@     q ~kOxq ~JQsq ~��w   ?@     q ~JFxq ~Z�sq ~��w   ?@     q ~Z�xq ~^sq ~��w   ?@     q ~^xq ~2{sq ~��w   ?@     q ~2pxq ~}-sq ~��w   ?@     q ~}"xq ~vsq ~��w   ?@     q ~u�xq ~_�sq ~��w   ?@     q ~_�xq ~RJsq ~��w   ?@     q ~R?xq ~C�sq ~��w   ?@     q ~C�xq ~��sq ~��w   ?@     q ~��xq ~p-sq ~��w   ?@     q ~p q ~��xq ~nwsq ~��w   ?@     q ~nixq ~�sq ~��w   ?@     q ~�xq ~@�sq ~��w   ?@     q ~@�xq ~�sq ~��w   ?@     q ~�xq ~Ovsq ~��w   ?@     q ~�\q ~Oixq ~(fsq ~��w   ?@     q ~(Yxq ~]sq ~��w   ?@     q ~Wxq ~c sq ~��w   ?@     q ~b�xq ~:�sq ~��w   ?@     q ~:�xq ~Zsq ~��w   ?@     q ~Zq ~'�xq ~J�sq ~��w   ?@     q ~J�xq ~;�sq ~��w   ?@     q ~;�xq ~nsq ~��w   ?@     q ~cxq ~Dlsq ~��w   ?@     q ~D^xq ~r&sq ~��w   ?@     q ~rxq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�xq ~tsq ~��w   ?@     q ~gq ~:dq ~C�xq ~{�sq ~��w   ?@     q ~{�q ~ �xq ~E�sq ~��w   ?@     q ~E�xq ~�>sq ~��w   ?@     q ~�3xq ~F�sq ~��w   ?@     q ~F�xq ~\sq ~��w   ?@     q ~\q ~l�xq ~0-sq ~��w   ?@     q ~0"xq ~9�sq ~��w   ?@     q ~9�xq ~sq ~��w   ?@     q ~�q ~C^xq ~Lsq ~��w   ?@     q ~Axq ~>$sq ~��w   ?@     q ~>xq ~v�sq ~��w   ?@     q ~v�xq ~k�sq ~��w   ?@     q ~k�xq ~{�sq ~��w   ?@     q ~{�xq ~@�sq ~��w   ?@     q ~@�xq ~/�sq ~��w   ?@     q ~/�xq ~��sq ~��w   ?@     q ~p�q ~��xq ~J�sq ~��w   ?@     q ~J�xq ~mpsq ~��w   ?@     q ~mexq ~]?sq ~��w   ?@     q ~]4xq ~��sq ~��w   ?@     q ~��q ~!xq ~�sq ~��w   ?@     q ~��q ~R�q ~9?q ~vq ~6xq ~vsq ~��w   ?@     q ~vxq ~n�sq ~��w   ?@     q ~n�xq ~8Fsq ~��w   ?@     q ~88xq ~_�sq ~��w   ?@     q ~_�xq ~Ywsq ~��w   ?@     q ~Ylxq ~�Vsq ~��w   ?@     q ~�Kxq ~ssq ~��w   ?@     q ~�q ~sxq ~�sq ~��w   ?@     q ~/gq ~�
xq ~
sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~_$sq ~��w   ?@     q ~_xq ~Psq ~��w   ?@     q ~Pxq ~xsq ~��w   ?@     q ~mxq ~j�sq ~��w   ?@     q ~j�xq ~s�sq ~��w   ?@     q ~s�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�q ~P_xq ~#asq ~��w   ?@     q ~#Vxq ~�sq ~��w   ?@     q ~�xq ~w	sq ~��w   ?@     q ~v�q ~K�xq ~{2sq ~��w   ?@     q ~{'q ~[xq ~wOsq ~��w   ?@     q ~wDq ~Uxq ~��sq ~��w   ?@     q ~��xq ~D�sq ~��w   ?@     q ~D�xq ~Ksq ~��w   ?@     q ~k�q ~=xq ~|sq ~��w   ?@     q ~{�xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�xq ~	qsq ~��w   ?@     q ~	cxq ~{�sq ~��w   ?@     q ~{�xq ~L�sq ~��w   ?@     q ~L�xq ~�,sq ~��w   ?@     q ~�!xq ~%-sq ~��w   ?@     q ~%"xq ~2�sq ~��w   ?@     q ~2}xq ~A�sq ~��w   ?@     q ~A�xq ~j�sq ~��w   ?@     q ~bq ~j�xq ~q�sq ~��w   ?@     q ~q�xq ~{sq ~��w   ?@     q ~{xq ~h�sq ~��w   ?@     q ~h�xq ~.�sq ~��w   ?@     q ~.�xq ~N�sq ~��w   ?@     q ~A�q ~N�xq ~insq ~��w   ?@     q ~i`q ~q4xq ~Nsq ~��w   ?@     q ~Nxq ~��sq ~��w   ?@     q ~��xq ~}�sq ~��w   ?@     q ~q ~}�xq ~\�sq ~��w   ?@     q ~\�xq ~t�sq ~��w   ?@     q ~t�xq ~R!sq ~��w   ?@     q ~Rq ~	�xq ~R�sq ~��w   ?@     q ~R�xq ~
>sq ~��w   ?@     q ~
0xq ~u�sq ~��w   ?@     q ~u�xq ~�sq ~��w   ?@     q ~�xq ~<�sq ~��w   ?@     q ~<�xq ~>vsq ~��w   ?@     q ~>pxq ~{�sq ~��w   ?@     q ~{�q ~*�xq ~msq ~��w   ?@     q ~�q ~l�xq ~25sq ~��w   ?@     q ~2'xq ~Dsq ~��w   ?@     q ~6xq ~V<sq ~��w   ?@     q ~V1xq ~�"sq ~��w   ?@     q ~�xq ~K sq ~��w   ?@     q ~J�xq ~i<sq ~��w   ?@     q ~i1xq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~Wsq ~��w   ?@     q ~�bq ~W xq ~G^sq ~��w   ?@     q ~�@q ~GSxq ~��sq ~��w   ?@     q ~��xq ~?wsq ~��w   ?@     q ~?lq ~xwxq ~mIsq ~��w   ?@     q ~m>xq ~m�sq ~��w   ?@     q ~m�xq ~3sq ~��w   ?@     q ~3xq ~��sq ~��w   ?@     q ~��xq ~9sq ~��w   ?@     q ~+xq ~�sq ~��w   ?@     q ~{xq ~L�sq ~��w   ?@     q ~L�q ~�)xq ~��sq ~��w   ?@     q ~D q ~��xq ~f�sq ~��w   ?@     q ~f�xq ~��sq ~��w   ?@     q ~��xq ~&�sq ~��w   ?@     q ~&�q ~DVxq ~-�sq ~��w   ?@     q ~-�xq ~X�sq ~��w   ?@     q ~X�xq ~�sq ~��w   ?@     q ~�
xq ~J�sq ~��w   ?@     q ~J�xq ~EFsq ~��w   ?@     q ~E@xq ~��sq ~��w   ?@     q ~��xq ~<�sq ~��w   ?@     q ~<�xq ~�asq ~��w   ?@     q ~�Vxq ~B�sq ~��w   ?@     q ~B�xq ~z�sq ~��w   ?@     q ~z�xq ~!Asq ~��w   ?@     q ~!3xq ~L0sq ~��w   ?@     q ~L%xq ~nKsq ~��w   ?@     q ~n@xq ~n1sq ~��w   ?@     q ~n&xq ~�9sq ~��w   ?@     q ~�q ~�.xq ~A�sq ~��w   ?@     q ~A�xq ~[}sq ~��w   ?@     q ~[rxq ~ �sq ~��w   ?@     q ~ |xq ~Isq ~��w   ?@     q ~Ixq ~e�sq ~��w   ?@     q ~ezxq ~;sq ~��w   ?@     q ~-q ~1�xq ~ <sq ~��w   ?@     q ~Yq ~ /xq ~�sq ~��w   ?@     q ~�xq ~e�sq ~��w   ?@     q ~e�xq ~;4sq ~��w   ?@     q ~�tq ~;'xq ~Ssq ~��w   ?@     q ~S xq ~=Gsq ~��w   ?@     q ~=<xq ~LWsq ~��w   ?@     q ~LLxq ~:�sq ~��w   ?@     q ~:�xq ~d�sq ~��w   ?@     q ~d�xq ~�>sq ~��w   ?@     q ~�3xq ~Hsq ~��w   ?@     q ~=xq ~d�sq ~��w   ?@     q ~d|xq ~$�sq ~��w   ?@     q ~$�xq ~sq ~��w   ?@     q ~xq ~qsq ~��w   ?@     q ~ixq ~�sq ~��w   ?@     q ~��xq ~\Ysq ~��w   ?@     q ~\Kxq ~�Nsq ~��w   ?@     q ~��q ~�Cxq ~|sq ~��w   ?@     q ~|xq ~H�sq ~��w   ?@     q ~I~q ~H�xq ~�sq ~��w   ?@     q ~�q ~; xq ~Y�sq ~��w   ?@     q ~+�q ~Y�q ~��xq ~Dsq ~��w   ?@     q ~�q ~Dxq ~w�sq ~��w   ?@     q ~w�xq ~��sq ~��w   ?@     q ~��xq ~f�sq ~��w   ?@     q ~�q ~f�xq ~sq ~��w   ?@     q ~��q ~�xq ~`gsq ~��w   ?@     q ~`\xq ~Lsq ~��w   ?@     q ~>xq ~&Qsq ~��w   ?@     q ~&Fxq ~\sq ~��w   ?@     q ~Nxq ~&7sq ~��w   ?@     q ~&,xq ~��sq ~��w   ?@     q ~��xq ~I�sq ~��w   ?@     q ~I�xq ~i{sq ~��w   ?@     q ~ipxq ~0�sq ~��w   ?@     q ~0zxq ~&�sq ~��w   ?@     q ~rq ~&�xq ~#qsq ~��w   ?@     q ~#cxq ~�usq ~��w   ?@     q ~�jxq ~�sq ~��w   ?@     q ~uxq ~�dsq ~��w   ?@     q ~�Yxq ~{�sq ~��w   ?@     q ~{�xq ~:Hsq ~��w   ?@     q ~:=xq ~q�sq ~��w   ?@     q ~q�xq ~� sq ~��w   ?@     q ~�xq ~@Nsq ~��w   ?@     q ~@Cxq ~sq ~��w   ?@     q ~qxq ~6esq ~��w   ?@     q ~6Zxq ~]sq ~��w   ?@     q ~��q ~]q ~q�xq ~��sq ~��w   ?@     q ~��xq ~_�sq ~��w   ?@     q ~_�xq ~Q.sq ~��w   ?@     q ~Q#xq ~R�sq ~��w   ?@     q ~R�xq ~K�sq ~��w   ?@     q ~K�xq ~sq ~��w   ?@     q ~xq ~x�sq ~��w   ?@     q ~x�q ~�xq ~.Esq ~��w   ?@     q ~apq ~.:xq ~k�sq ~��w   ?@     q ~k�xq ~-Wsq ~��w   ?@     q ~-Ixq ~)Ksq ~��w   ?@     q ~)@xq ~sq ~��w   ?@     q ~xq ~s�sq ~��w   ?@     q ~s�xq ~b�sq ~��w   ?@     q ~bvxq ~
�sq ~��w   ?@     q ~
�xq ~�sq ~��w   ?@     q ~��q ~p�xq ~p�sq ~��w   ?@     q ~p�q ~(Ixq ~{�sq ~��w   ?@     q ~{�xq ~�sq ~��w   ?@     q ~�xq ~Msq ~��w   ?@     q ~Mxq ~F:sq ~��w   ?@     q ~F/xq ~5Osq ~��w   ?@     q ~5Dxq ~V�sq ~��w   ?@     q ~Vwxq ~i�sq ~��w   ?@     q ~i�xq ~lWsq ~��w   ?@     q ~[eq ~lIxq ~e�sq ~��w   ?@     q ~e�xq ~p�sq ~��w   ?@     q ~p�xq ~Adsq ~��w   ?@     q ~AYxq ~��sq ~��w   ?@     q ~��xq ~uysq ~��w   ?@     q ~unxq ~t'sq ~��w   ?@     q ~txq ~k
sq ~��w   ?@     q ~Qq ~j�xq ~isq ~��w   ?@     q ~ "q ~h�xq ~Q�sq ~��w   ?@     q ~Q�q ~,ixq ~�;sq ~��w   ?@     q ~�0xq ~3�sq ~��w   ?@     q ~3�xq ~V�sq ~��w   ?@     q ~V�xq ~Dsq ~��w   ?@     q ~6xq ~�sq ~��w   ?@     q ~�xq ~~sq ~��w   ?@     q ~~xq ~j�sq ~��w   ?@     q ~j�xq ~Asq ~��w   ?@     q ~�;q ~Axq ~E�sq ~��w   ?@     q ~E�xq ~m�sq ~��w   ?@     q ~m�xq ~N�sq ~��w   ?@     q ~N�xq ~�sq ~��w   ?@     q ~�xq ~X�sq ~��w   ?@     q ~X�q ~q�xq ~jsq ~��w   ?@     q ~jq ~V�xq ~+1sq ~��w   ?@     q ~+&xq ~��sq ~��w   ?@     q ~��q ~�xq ~?�sq ~��w   ?@     q ~?�xq ~9=sq ~��w   ?@     q ~92xq ~Psq ~��w   ?@     q ~Pxq ~�sq ~��w   ?@     q ~�xq ~U,sq ~��w   ?@     q ~Uq ~'xq ~T�sq ~��w   ?@     q ~Txq ~Z�sq ~��w   ?@     q ~Z�xq ~�sq ~��w   ?@     q ~|xq ~4sq ~��w   ?@     q ~4xq ~2�sq ~��w   ?@     q ~2�xq ~w�sq ~��w   ?@     q ~w�xq ~�Usq ~��w   ?@     q ~�Jxq ~u�sq ~��w   ?@     q ~-q ~t�q ~q ~s,q ~u�xq ~{�sq ~��w   ?@     q ~Fcq ~{�xq ~@�sq ~��w   ?@     q ~@�q ~O@xq ~WLsq ~��w   ?@     q ~WAxq ~
qsq ~��w   ?@     q ~
cxq ~G�sq ~��w   ?@     q ~G�xq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~t�sq ~��w   ?@     q ~t�xq ~ �sq ~��w   ?@     q ~ �xq ~lsq ~��w   ?@     q ~vq ~^xq ~Qsq ~��w   ?@     q ~Cxq ~P�sq ~��w   ?@     q ~P�xq ~tsq ~��w   ?@     q ~V�q ~t q ~�xq ~�sq ~��w   ?@     q ~�xq ~%sq ~��w   ?@     q ~%xq ~sq ~��w   ?@     q ~ xq ~n\sq ~��w   ?@     q ~nNxq ~4�sq ~��w   ?@     q ~4�xq ~%�sq ~��w   ?@     q ~%�xq ~6Hsq ~��w   ?@     q ~6=xq ~�sq ~��w   ?@     q ~�xq ~i�sq ~��w   ?@     q ~i�xq ~psq ~��w   ?@     q ~yq ~pxq ~*�sq ~��w   ?@     q ~*�xq ~�:sq ~��w   ?@     q ~�/xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~�q ~@�xq ~fWsq ~��w   ?@     q ~)�q ~fIxq ~S�sq ~��w   ?@     q ~S�xq ~m<sq ~��w   ?@     q ~m1xq ~p�sq ~��w   ?@     q ~p�xq ~�sq ~��w   ?@     q ~{xq ~PPsq ~��w   ?@     q ~PExq ~K6sq ~��w   ?@     q ~K)q ~@�xq ~8�sq ~��w   ?@     q ~8�xq ~w�sq ~��w   ?@     q ~w�xq ~<sq ~��w   ?@     q ~<
xq ~O�sq ~��w   ?@     q ~��q ~Oxxq ~<�sq ~��w   ?@     q ~<�xq ~esq ~��w   ?@     q ~Wq ~<�xq ~sq ~��w   ?@     q ~~�xq ~&sq ~��w   ?@     q ~}�q ~&xq ~Aqsq ~��w   ?@     q ~Afxq ~s�sq ~��w   ?@     q ~s�xq ~~�sq ~��w   ?@     q ~~uxq ~f�sq ~��w   ?@     q ~f�xq ~U
sq ~��w   ?@     q ~T�xq ~e<sq ~��w   ?@     q ~e/q ~?xq ~Dsq ~��w   ?@     q ~Qq ~5xq ~n�sq ~��w   ?@     q ~n�xq ~D�sq ~��w   ?@     q ~D�xq ~Fsq ~��w   ?@     q ~8xq ~nsq ~��w   ?@     q ~cq ~Bxq ~sq ~��w   ?@     q ~/�q ~ xq ~:sq ~��w   ?@     q ~,xq ~K�sq ~��w   ?@     q ~K�xq ~D�sq ~��w   ?@     q ~D�xq ~7Wsq ~��w   ?@     q ~Uq ~7Lxq ~]%sq ~��w   ?@     q ~]xq ~_�sq ~��w   ?@     q ~_�q ~�xq ~�sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~wq ~�uxq ~BPsq ~��w   ?@     q ~BExq ~Y�sq ~��w   ?@     q ~-�q ~Y�xq ~MWsq ~��w   ?@     q ~MIxq ~s\sq ~��w   ?@     q ~sQxq ~.�sq ~��w   ?@     q ~.�xq ~�Msq ~��w   ?@     q ~)�q ~�@xq ~�sq ~��w   ?@     q ~�xq ~W�sq ~��w   ?@     q ~W�xq ~7�sq ~��w   ?@     q ~7�xq ~�sq ~��w   ?@     q ~@&q ~�xq ~}�sq ~��w   ?@     q ~}�q ~|xq ~��sq ~��w   ?@     q ~��xq ~e-sq ~��w   ?@     q ~e"xq ~�sq ~��w   ?@     q ~�xq ~?�sq ~��w   ?@     q ~?�xq ~S�sq ~��w   ?@     q ~S�xq ~��sq ~��w   ?@     q ~��q ~XRxq ~:�sq ~��w   ?@     q ~:�xq ~n�sq ~��w   ?@     q ~nzq ~q�xq ~sq ~��w   ?@     q ~xq ~�{sq ~��w   ?@     q ~�sxq ~COsq ~��w   ?@     q ~CDxq ~�sq ~��w   ?@     q ~�$q ~�xq ~U�sq ~��w   ?@     q ~U�xq ~u5sq ~��w   ?@     q ~u*xq ~fGsq ~��w   ?@     q ~f<xq ~�Osq ~��w   ?@     q ~�Dxq ~gsq ~��w   ?@     q ~gxq ~W2sq ~��w   ?@     q ~W'xq ~xYsq ~��w   ?@     q ~xKq ~%xq ~�\sq ~��w   ?@     q ~�Qxq ~�"sq ~��w   ?@     q ~U;q ~�xq ~"�sq ~��w   ?@     q ~"�xq ~|sq ~��w   ?@     q ~|q ~�3xq ~L�sq ~��w   ?@     q ~�q ~L�xq ~Csq ~��w   ?@     q ~C	xq ~dsq ~��w   ?@     q ~Yxq ~6�sq ~��w   ?@     q ~6�xq ~"6sq ~��w   ?@     q ~"(xq ~�qsq ~��w   ?@     q ~�fxq ~`%sq ~��w   ?@     q ~`xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~$�q ~zxq ~�tsq ~��w   ?@     q ~�fq ~L�xq ~5'sq ~��w   ?@     q ~5xq ~��sq ~��w   ?@     q ~��xq ~4sq ~��w   ?@     q ~4txq ~A~sq ~��w   ?@     q ~Asxq ~T�sq ~��w   ?@     q ~d<q ~T�xq ~b-sq ~��w   ?@     q ~b"xq ~5\sq ~��w   ?@     q ~5Qq ~�9xq ~(sq ~��w   ?@     q ~(xq ~!�sq ~��w   ?@     q ~8�q ~!�xq ~%�sq ~��w   ?@     q ~%�xq ~��sq ~��w   ?@     q ~l�q ~��xq ~�Gsq ~��w   ?@     q ~1�q ~�<xq ~(�sq ~��w   ?@     q ~(�xq ~C�sq ~��w   ?@     q ~C�xq ~>�sq ~��w   ?@     q ~>�xq ~"Vsq ~��w   ?@     q ~<eq ~"Hxq ~k�sq ~��w   ?@     q ~k�xq ~jlsq ~��w   ?@     q ~jaxq ~@�sq ~��w   ?@     q ~@�xq ~;�sq ~��w   ?@     q ~;�xq ~Vhsq ~��w   ?@     q ~?�q ~V]xq ~ozsq ~��w   ?@     q ~ooxq ~7gsq ~��w   ?@     q ~7Yxq ~4sq ~��w   ?@     q ~&xq ~Lsq ~��w   ?@     q ~L	q ~}/xq ~Gxsq ~��w   ?@     q ~Gmxq ~4sq ~��w   ?@     q ~'xq ~.sq ~��w   ?@     q ~�q ~.q ~\(xq ~^Isq ~��w   ?@     q ~^<q ~Vxq ~esq ~��w   ?@     q ~Wxq ~2sq ~��w   ?@     q ~2xq ~r�sq ~��w   ?@     q ~r�xq ~6,sq ~��w   ?@     q ~�q ~6xq ~y�sq ~��w   ?@     q ~y�xq ~rBsq ~��w   ?@     q ~r7xq ~�Hsq ~��w   ?@     q ~�=xq ~?Ysq ~��w   ?@     q ~?Qxq ~Csq ~��w   ?@     q ~5xq ~*�sq ~��w   ?@     q ~*�xq ~�sq ~��w   ?@     q ~�xq ~ sq ~��w   ?@     q ~xq ~#sq ~��w   ?@     q ~xq ~z�sq ~��w   ?@     q ~�q ~z�xq ~+�sq ~��w   ?@     q ~+�q ~	�xq ~#sq ~��w   ?@     q ~xq ~+sq ~��w   ?@     q ~+xq ~E�sq ~��w   ?@     q ~E�q ~<>xq ~) sq ~��w   ?@     q ~)xq ~�sq ~��w   ?@     q ~�xq ~sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~:sq ~��w   ?@     q ~,xq ~:�sq ~��w   ?@     q ~:�xq ~)sq ~��w   ?@     q ~)xq ~��sq ~��w   ?@     q ~��xq ~�sq ~��w   ?@     q ~4q ~�xq ~b�sq ~��w   ?@     q ~b�xq ~H�sq ~��w   ?@     q ~Q=q ~H�xq ~Fsq ~��w   ?@     q ~Fq ~
xq ~#�sq ~��w   ?@     q ~#�xq ~5�sq ~��w   ?@     q ~5�xq ~bsq ~��w   ?@     q ~a�xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~"~q ~A�q ~�xq ~*�sq ~��w   ?@     q ~*{xq ~;{sq ~��w   ?@     q ~;pxq ~)-sq ~��w   ?@     q ~)"xq ~C�sq ~��w   ?@     q ~Cxxq ~ sq ~��w   ?@     q ~xq ~K�sq ~��w   ?@     q ~Kyxq ~|�sq ~��w   ?@     q ~�q ~|�xq ~5�sq ~��w   ?@     q ~5�xq ~-�sq ~��w   ?@     q ~-�xq ~-7sq ~��w   ?@     q ~-,xq ~ansq ~��w   ?@     q ~wq ~aaxq ~�sq ~��w   ?@     q ~�xq ~9�sq ~��w   ?@     q ~9�xq ~ssq ~��w   ?@     q ~hxq ~b�sq ~��w   ?@     q ~b�xq ~Ssq ~��w   ?@     q ~Exq ~g&sq ~��w   ?@     q ~gxq ~	�sq ~��w   ?@     q ~	�xq ~XPsq ~��w   ?@     q ~XExq ~Ogsq ~��w   ?@     q ~O\xq ~vhsq ~��w   ?@     q ~v]xq ~6sq ~��w   ?@     q ~;�q ~-�q ~+q ~xq ~%�sq ~��w   ?@     q ~%�xq ~SLsq ~��w   ?@     q ~SAxq ~z�sq ~��w   ?@     q ~�/q ~z�xq ~Jusq ~��w   ?@     q ~Joxq ~Jsq ~��w   ?@     q ~Jxq ~�sq ~��w   ?@     q ~�xq ~ulsq ~��w   ?@     q ~uaxq ~,Zsq ~��w   ?@     q ~,Oq ~D�q ~j�xq ~5�sq ~��w   ?@     q ~5�xq ~O�sq ~��w   ?@     q ~O�q ~��q ~�xq ~Bsq ~��w   ?@     q ~4xq ~+$sq ~��w   ?@     q ~M�q ~i�q ~b�q ~+q ~�xq ~sq ~��w   ?@     q ~�q ~w(xq ~U�sq ~��w   ?@     q ~U�xq ~2sq ~��w   ?@     q ~Y�q ~$xq ~o�sq ~��w   ?@     q ~o�q ~%/xq ~k�sq ~��w   ?@     q ~k�xq ~w�sq ~��w   ?@     q ~w�q ~~�xq ~\sq ~��w   ?@     q ~Nq ~b>xq ~p:sq ~��w   ?@     q ~p/xq ~��sq ~��w   ?@     q ~��xq ~�]sq ~��w   ?@     q ~�Rxq ~hsq ~��w   ?@     q ~hxq ~pWsq ~��w   ?@     q ~��q ~pLxq ~P�sq ~��w   ?@     q ~?�q ~P�xq ~;asq ~��w   ?@     q ~;Vq ~pxq ~�sq ~��w   ?@     q ~�xq ~-�sq ~��w   ?@     q ~Suq ~-�xq ~�sq ~��w   ?@     q ~�xq ~I�sq ~��w   ?@     q ~I�xq ~P�sq ~��w   ?@     q ~P�q ~YRxq ~!Qsq ~��w   ?@     q ~!Dxq ~��sq ~��w   ?@     q ~��xq ~)�sq ~��w   ?@     q ~)�xq ~i�sq ~��w   ?@     q ~i�q ~E�xq ~O!sq ~��w   ?@     q ~Oxq ~@$sq ~��w   ?@     q ~@q ~#xq ~i^sq ~��w   ?@     q ~iSxq ~,sq ~��w   ?@     q ~!xq ~Csq ~��w   ?@     q ~B�xq ~%wsq ~��w   ?@     q ~%jxq ~	�sq ~��w   ?@     q ~	�xq ~7sq ~��w   ?@     q ~7xq ~!~sq ~��w   ?@     q ~!pxq ~Lsq ~��w   ?@     q ~>xq ~#Tsq ~��w   ?@     q ~#Ixq ~U�sq ~��w   ?@     q ~U�xq ~�ssq ~��w   ?@     q ~�hxq ~��sq ~��w   ?@     q ~��xq ~>�sq ~��w   ?@     q ~>�q ~�<q ~xq ~]
sq ~��w   ?@     q ~\�q ~y�xq ~4�sq ~��w   ?@     q ~4�xq ~t�sq ~��w   ?@     q ~t�xq ~�!sq ~��w   ?@     q ~�xq ~��sq ~��w   ?@     q ~��xq ~W�sq ~��w   ?@     q ~W�xq ~ �sq ~��w   ?@     q ~ �xq ~�sq ~��w   ?@     q ~��xq ~$?sq ~��w   ?@     q ~$1xq ~{|sq ~��w   ?@     q ~{qxq ~vsq ~��w   ?@     q ~vxq ~csq ~��w   ?@     q ~Xxq ~L=sq ~��w   ?@     q ~L2xq ~��sq ~��w   ?@     q ~�yq ~�Ixq ~p�sq ~��w   ?@     q ~psq ~�xq ~Hlsq ~��w   ?@     q ~Hfxq ~>�sq ~��w   ?@     q ~>�xq ~�sq ~��w   ?@     q ~zxq ~FTsq ~��w   ?@     q ~FIq ~��xq ~a�sq ~��w   ?@     q ~a�xq ~�sq ~��w   ?@     q ~zxq ~O�sq ~��w   ?@     q ~O�q ~D�xq ~%�sq ~��w   ?@     q ~%�xq ~�Tsq ~��w   ?@     q ~�Ixq ~/�sq ~��w   ?@     q ~/�xq ~_sq ~��w   ?@     q ~Txq ~jsq ~��w   ?@     q ~jq ~��xq ~<�sq ~��w   ?@     q ~q ~<�xq ~ysq ~��w   ?@     q ~nxq ~<�sq ~��w   ?@     q ~<uxq ~\sq ~��w   ?@     q ~\xq ~l�sq ~��w   ?@     q ~Dq ~lwxq ~Qesq ~��w   ?@     q ~QWxq ~"^sq ~��w   ?@     q ~"Xxq ~�sq ~��w   ?@     q ~�xq ~Asq ~��w   ?@     q ~2�q ~Axq ~.8sq ~��w   ?@     q ~.+q ~S�xq ~|Xsq ~��w   ?@     q ~|Jxq ~�;sq ~��w   ?@     q ~�0xq ~>sq ~��w   ?@     q ~=�xq ~!�sq ~��w   ?@     q ~!�xq ~,�sq ~��w   ?@     q ~,�xq ~t�sq ~��w   ?@     q ~t�xq ~Bsq ~��w   ?@     q ~A�xq ~usq ~��w   ?@     q ~gxq ~l�sq ~��w   ?@     q ~l�q ~zxq ~�sq ~��w   ?@     q ~�xq ~sq ~��w   ?@     q ~ �xq ~|�sq ~��w   ?@     q ~|�xq ~?5sq ~��w   ?@     q ~?*xq ~Csq ~��w   ?@     q ~8xq ~(Gsq ~��w   ?@     q ~(<xq ~|�sq ~��w   ?@     q ~|�xq ~r�sq ~��w   ?@     q ~r�xq ~��sq ~��w   ?@     q ~��xq ~sq ~��w   ?@     q ~xq ~j�sq ~��w   ?@     q ~j�xq ~�Osq ~��w   ?@     q ~�Dxq ~�sq ~��w   ?@     q ~�q ~�^xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�xq ~�Csq ~��w   ?@     q ~�8xq ~Xwsq ~��w   ?@     q ~Xlxq ~Ssq ~��w   ?@     q ~Sxq ~:|sq ~��w   ?@     q ~:qxq ~4Xsq ~��w   ?@     q ~4Mq ~P+q ~,@xq ~�sq ~��w   ?@     q ~�xq ~�|sq ~��w   ?@     q ~�qq ~_xq ~mcsq ~��w   ?@     q ~mXq ~�xq ~i�sq ~��w   ?@     q ~i�xq ~2�sq ~��w   ?@     q ~2�xq ~Zlsq ~��w   ?@     q ~Zaxq ~e�sq ~��w   ?@     q ~e�xq ~j,sq ~��w   ?@     q ~j!xq ~`�sq ~��w   ?@     q ~`�xq ~v�sq ~��w   ?@     q ~v�xq ~]sq ~��w   ?@     q ~Oxq ~.�sq ~��w   ?@     q ~.�xq ~sq ~��w   ?@     q ~	xq ~f:sq ~��w   ?@     q ~Y�q ~f/xq ~ysq ~��w   ?@     q ~yxq ~@�sq ~��w   ?@     q ~@�xq ~P�sq ~��w   ?@     q ~P�xq ~7�sq ~��w   ?@     q ~7�xq ~Z�sq ~��w   ?@     q ~Z�xq ~7Isq ~��w   ?@     q ~7;xq ~tsq ~��w   ?@     q ~ttxq ~}�sq ~��w   ?@     q ~}�xq ~�sq ~��w   ?@     q ~�xq ~Q�sq ~��w   ?@     q ~Q�xq ~2sq ~��w   ?@     q ~$xq ~>sq ~��w   ?@     q ~>xq ~5	sq ~��w   ?@     q ~B_q ~�q ~�lq ~jRq ~4�xq ~V�sq ~��w   ?@     q ~V�xq ~d�sq ~��w   ?@     q ~d�xq ~c,sq ~��w   ?@     q ~cxq ~n
sq ~��w   ?@     q ~m�xq ~2�sq ~��w   ?@     q ~2�xq ~F,sq ~��w   ?@     q ~Fq ~�xq ~e�sq ~��w   ?@     q ~e�xq ~`�sq ~��w   ?@     q ~`�q ~@Pxq ~2asq ~��w   ?@     q ~2Vxq ~w�sq ~��w   ?@     q ~w�q ~�Jxq ~�sq ~��w   ?@     q ~�xq ~P�sq ~��w   ?@     q ~P�xq ~u�sq ~��w   ?@     q ~u�q ~]Axq ~B5sq ~��w   ?@     q ~B/xq ~o]sq ~��w   ?@     q ~e�q ~oRxq ~ sq ~��w   ?@     q ~�xq ~o(sq ~��w   ?@     q ~o xq ~�sq ~��w   ?@     q ~xxq ~5ysq ~��w   ?@     q ~5nxq ~�sq ~��w   ?@     q ~��xq ~k�sq ~��w   ?@     q ~k�xq ~Lsq ~��w   ?@     q ~>q ~\hxq ~eLsq ~��w   ?@     q ~e>xq ~`sq ~��w   ?@     q ~Uxq ~)Usq ~��w   ?@     q ~)Mxq ~�sq ~��w   ?@     q ~�xq ~7�sq ~��w   ?@     q ~7�xq ~6sq ~��w   ?@     q ~�_q ~6xq ~l(sq ~��w   ?@     q ~lxq ~I�sq ~��w   ?@     q ~I�xq ~6sq ~��w   ?@     q ~6xq ~Z�sq ~��w   ?@     q ~Z{xq ~��sq ~��w   ?@     q ~��xq ~|�sq ~��w   ?@     q ~|�xq ~Jmsq ~��w   ?@     q ~Jbxq ~0sq ~��w   ?@     q ~aq ~��q ~%q ~G�xq ~��sq ~��w   ?@     q ~��xq ~(�sq ~��w   ?@     q ~(�xq ~��sq ~��w   ?@     q ~��xq ~U�sq ~��w   ?@     q ~U�xq ~vsq ~��w   ?@     q ~kxq ~�sq ~��w   ?@     q ~g�q ~�xq ~$�sq ~��w   ?@     q ~$�q ~"�xq ~��sq ~��w   ?@     q ~��xq ~osq ~��w   ?@     q ~oxq ~Osq ~��w   ?@     q ~O	xq ~e�sq ~��w   ?@     q ~e�xq ~��sq ~��w   ?@     q ~��xq ~_|sq ~��w   ?@     q ~_qxq ~�(sq ~��w   ?@     q ~�xq ~sq ~��w   ?@     q ~�q ~i�xq ~=�sq ~��w   ?@     q ~=�xq ~��sq ~��w   ?@     q ~��xq ~  sq ~��w   ?@     q ~�q ~ xq ~D�sq ~��w   ?@     q ~D�xq ~m}sq ~��w   ?@     q ~mrxq ~��sq ~��w   ?@     q ~��xq ~�Hsq ~��w   ?@     q ~�=xq ~%hsq ~��w   ?@     q ~%]xq ~=dsq ~��w   ?@     q ~=Yxq ~;�sq ~��w   ?@     q ~;�xq ~Z�sq ~��w   ?@     q ~Z�xq ~=:sq ~��w   ?@     q ~I)q ~=-xq ~.�sq ~��w   ?@     q ~.rxq ~}Wsq ~��w   ?@     q ~}Iq ~Pxq ~0sq ~��w   ?@     q ~/�xq ~��sq ~��w   ?@     q ~��q ~=nxq ~��sq ~��w   ?@     q ~�~xq ~Upsq ~��w   ?@     q ~Uexq ~O�sq ~��w   ?@     q ~O�q ~�xq ~i/sq ~��w   ?@     q ~i$xq ~�sq ~��w   ?@     q ~�xq ~�sq ~��w   ?@     q ~�q ~��xq ~lsq ~��w   ?@     q ~`�q ~lxq ~Y�sq ~��w   ?@     q ~Y�xq ~_>sq ~��w   ?@     q ~_3xq ~\�sq ~��w   ?@     q ~\�xq ~N�sq ~��w   ?@     q ~N�q ~T�xq ~g�sq ~��w   ?@     q ~g�xq ~-sq ~��w   ?@     q ~�Rq ~-xq ~4Ksq ~��w   ?@     q ~V�q ~4>xq ~&�sq ~��w   ?@     q ~&�xq ~^�sq ~��w   ?@     q ~^sxq ~4�sq ~��w   ?@     q ~4�xq ~sq ~��w   ?@     q ~xq ~wBsq ~��w   ?@     q ~w7xq ~y�sq ~��w   ?@     q ~~4q ~y�xq ~3�sq ~��w   ?@     q ~3�xq ~��sq ~��w   ?@     q ~��xq ~6�sq ~��w   ?@     q ~6�xq ~Z_sq ~��w   ?@     q ~ZTxq ~H0sq ~��w   ?@     q ~H%xq ~dQsq ~��w   ?@     q ~dFxq ~3�sq ~��w   ?@     q ~3�xq ~j{sq ~��w   ?@     q ~jnq ~��xq ~|�sq ~��w   ?@     q ~|�xq ~G�sq ~��w   ?@     q ~41q ~G�xq ~�sq ~��w   ?@     q ~�q ~x/xq ~sq ~��w   ?@     q ~l�q ~xq ~X�sq ~��w   ?@     q ~X�xq ~<�sq ~��w   ?@     q ~<�xq ~�sq ~��w   ?@     q ~�xq ~7�sq ~��w   ?@     q ~7�xq ~\�sq ~��w   ?@     q ~\�xq ~��sq ~��w   ?@     q ~��xq ~N<sq ~��w   ?@     q ~N1xq ~tsq ~��w   ?@     q ~ixq ~/=sq ~��w   ?@     q ~//xq ~<<sq ~��w   ?@     q ~<1xq ~�sq ~��w   ?@     q ~�q ~M�xq ~�bsq ~��w   ?@     q ~�Wxq ~iQsq ~��w   ?@     q ~iFxq ~�sq ~��w   ?@     q ~�xq ~OZsq ~��w   ?@     q ~OOxq ~N�sq ~��w   ?@     q ~N�xq ~�sq ~��w   ?@     q ~�xq ~fsq ~��w   ?@     q ~e�xq ~7�sq ~��w   ?@     q ~7�xq ~�sq ~��w   ?@     q ~�xq ~K'sq ~��w   ?@     q ~Kxq ~-*sq ~��w   ?@     q ~-xq ~zIsq ~��w   ?@     q ~z>xq ~��sq ~��w   ?@     q ~��xq ~Bwsq ~��w   ?@     q ~Biq ~�xq ~3�sq ~��w   ?@     q ~3�xq ~Gksq ~��w   ?@     q ~G`xq ~Vusq ~��w   ?@     q ~q ~Vjxq ~sq ~��w   ?@     q ~xq ~��sq ~��w   ?@     q ~��xq ~@Asq ~��w   ?@     q ~@6xq ~�ysq ~��w   ?@     q ~�nxq ~�sq ~��w   ?@     q ~�
xq ~Fsq ~��w   ?@     q ~E�xq ~yisq ~��w   ?@     q ~y^xq ~r�sq ~��w   ?@     q ~r�xq ~^�sq ~��w   ?@     q ~^�xq ~ �sq ~��w   ?@     q ~ �q ~KExq ~:.sq ~��w   ?@     q ~:#q ~�xq ~r�sq ~��w   ?@     q ~r�xq ~/sq ~��w   ?@     q ~!xq ~\�sq ~��w   ?@     q ~=q ~\�xq ~��sq ~��w   ?@     q ~��q ~8xq ~�sq ~��w   ?@     q ~�xq ~P�sq ~��w   ?@     q ~P�xq ~�Wsq ~��w   ?@     q ~wq ~�Jxq ~~fsq ~��w   ?@     q ~~[xq ~\�sq ~��w   ?@     q ~\�xq ~3^sq ~��w   ?@     q ~3Sxq ~Z4sq ~��w   ?@     q ~Z,xq ~`sq ~��w   ?@     q ~I�q ~_�q ~Lfxq ~)�sq ~��w   ?@     q ~q ~)�q ~��xq ~o�sq ~��w   ?@     q ~o�xq ~DTsq ~��w   ?@     q ~DIxq ~�sq ~��w   ?@     q ~	�q ~�xq ~b�sq ~��w   ?@     q ~�q ~b�xq ~HWsq ~��w   ?@     q ~HLxq ~0=sq ~��w   ?@     q ~0/xq ~	�sq ~��w   ?@     q ~	�q ~h�xq ~Esq ~��w   ?@     q ~Exq ~(:sq ~��w   ?@     q ~(/xq ~n�sq ~��w   ?@     q ~n�xq ~�'sq ~��w   ?@     q ~g(q ~�xq ~Ksq ~��w   ?@     q ~Kxq ~LJsq ~��w   ?@     q ~zq ~L?xq ~�sq ~��w   ?@     q ~�xq ~$�sq ~��w   ?@     q ~$�q ~�rxq ~�sq ~��w   ?@     q ~�xq ~�hsq ~��w   ?@     q ~�]xq ~c�sq ~��w   ?@     q ~c�xq ~~�sq ~��w   ?@     q ~m�q ~~�xq ~FGsq ~��w   ?@     q ~F<xq ~q�sq ~��w   ?@     q ~quq ~U�xq ~�sq ~��w   ?@     q ~vxq ~�sq ~��w   ?@     q ~c�q ~�xq ~vKsq ~��w   ?@     q ~v@xq ~i�sq ~��w   ?@     q ~i�xq ~X�sq ~��w   ?@     q ~X�xq ~Usq ~��w   ?@     q ~Gxq ~k@sq ~��w   ?@     q ~k5xq ~�sq ~��w   ?@     q ~�q ~.�xq ~Xjsq ~��w   ?@     q ~X_xq ~Osq ~��w   ?@     q ~Bxq ~\Hsq ~��w   ?@     q ~\Bxq ~2�sq ~��w   ?@     q ~2�xq ~F�sq ~��w   ?@     q ~F�xq ~�sq ~��w   ?@     q ~�xq ~`�sq ~��w   ?@     q ~`�xq ~�sq ~��w   ?@     q ~xxq ~]�sq ~��w   ?@     q ~]�xq ~	sq ~��w   ?@     q ~�xxsq ~ C?@     w       q ~u�sq ~��w   ?@     q ~B�q ~]�q ~�q ~��q ~u�xq ~��sq ~��w   @?@     &q ~��q ~q�q ~~!q ~_q ~L�q ~|�q ~~�q ~F�q ~q ~eq ~M�q ~. q ~|~q ~+q ~Eq ~��q ~X;q ~$q ~UZq ~O�q ~�wq ~�q ~raq ~7jq ~��q ~K�q ~Suq ~i�q ~=�q ~s,q ~1q ~��q ~q ~nq ~oq ~Vq ~0q ~p�xq ~M�sq ~��w   ?@     q ~M�q ~+q ~DVxq ~@�sq ~��w   �?@     Tq ~+�q ~��q ~tq ~X�q ~T�q ~0�q ~�q ~|uq ~>�q ~n�q ~d�q ~��q ~�Oq ~��q ~�yq ~0�q ~~�q ~*�q ~Xyq ~>pq ~p�q ~;�q ~@�q ~\Bq ~@�q ~aq ~z�q ~�q ~Hfq ~Joq ~��q ~Q�q ~"�q ~i�q ~xq ~qq ~-�q ~x�q ~q ~V�q ~��q ~R�q ~Q�q ~V�q ~E@q ~6�q ~{Aq ~q ~�q ~Hnq ~n@q ~Xq ~x�q ~*�q ~s�q ~�q ~t�q ~"Xq ~2�q ~�Dq ~q ~^q ~<>q ~{q ~!�q ~Fq ~�q ~-�q ~7q ~e�q ~2�q ~	�q ~_�q ~Wq ~0�q ~��q ~Uq ~Qq ~B/q ~�Cq ~^Xq ~O�q ~d'q ~o|xq ~1zsq ~��w   ?@    	[q ~L	q ~�q ~D�q ~M�q ~Xq ~t�q ~Yyq ~�q ~i�q ~^�q ~1&q ~�<q ~R�q ~:�q ~c<q ~D�q ~Q�q ~j�q ~(�q ~�Vq ~Z7q ~8�q ~=}q ~d�q ~vq ~Y�q ~��q ~_&q ~l�q ~f�q ~j�q ~�q ~z>q ~/Mq ~	�q ~]�q ~�3q ~K�q ~~4q ~o�q ~�9q ~�q ~�q ~[�q ~D q ~|�q ~J�q ~!�q ~/?q ~j�q ~2Eq ~r�q ~2}q ~�q ~e\q ~q ~n3q ~~�q ~f�q ~�q ~3q ~mKq ~I�q ~sq ~`�q ~\(q ~yq ~a�q ~�q ~z�q ~3,q ~�q ~�q ~!�q ~��q ~��q ~N�q ~Eq ~o�q ~IPq ~ceq ~\�q ~[q ~	cq ~�Jq ~6.q ~4>q ~��q ~(�q ~T,q ~i}q ~�@q ~7tq ~p�q ~}�q ~r(q ~.rq ~Znq ~ q ~Plq ~q ~��q ~L�q ~q ~;}q ~k�q ~�0q ~_�q ~#�q ~9�q ~41q ~;Vq ~Y�q ~��q ~^q ~�q ~�Mq ~6�q ~�q ~A�q ~q ~*�q ~+�q ~q ~+~q ~=�q ~�q ~X,q ~��q ~92q ~Vq ~@lq ~�q ~"�q ~I�q ~Ylq ~P�q ~niq ~Z{q ~,q ~q4q ~�q ~�q ~qhq ~4q ~6tq ~O�q ~q ~Wq ~��q ~:�q ~c�q ~��q ~�fq ~5q ~Jq ~;�q ~g�q ~8Yq ~fYq ~:Wq ~u�q ~8Hq ~n�q ~k�q ~5Qq ~q ~9�q ~x[q ~�Xq ~K�q ~!q ~�lq ~e/q ~_qq ~q�q ~skq ~��q ~F�q ~O\q ~��q ~+�q ~��q ~�q ~f�q ~{Wq ~3�q ~}q ~k�q ~8�q ~A�q ~!3q ~Yq ~!�q ~uDq ~p�q ~a�q ~`vq ~;�q ~F�q ~giq ~Vq ~pLq ~F�q ~2�q ~m�q ~��q ~��q ~V�q ~iq ~�q ~uq ~0"q ~EIq ~1�q ~2�q ~��q ~�3q ~&�q ~nq ~;q ~,q ~q�q ~)Xq ~c�q ~�q ~O�q ~+Pq ~K�q ~�q ~v q ~Dyq ~-,q ~��q ~)�q ~J�q ~X�q ~\q ~5nq ~-q ~l�q ~1�q ~P�q ~r�q ~3}q ~LYq ~s4q ~=-q ~F�q ~6�q ~b/q ~�=q ~�q ~@	q ~7.q ~q ~ q ~DIq ~k(q ~$jq ~B�q ~S�q ~x�q ~G�q ~�q ~G�q ~N�q ~;�q ~]�q ~%�q ~��q ~1rq ~HYq ~��q ~q ~Ckq ~#�q ~�eq ~�@q ~q ~E�q ~9Yq ~\uq ~xq ~mq ~3�q ~E�q ~�Uq ~Y8q ~[Xq ~T<q ~>�q ~q�q ~�nq ~�q ~q�q ~o�q ~q ~�q ~!pq ~-q ~�q ~�q ~C�q ~d�q ~��q ~$�q ~d�q ~{q ~/�q ~Pq ~${q ~^"q ~zq ~Zq ~q ~Tq ~��q ~{�q ~�q ~,�q ~�q ~X q ~k�q ~kBq ~�0q ~�q ~��q ~m�q ~2cq ~tKq ~�q ~^fq ~LLq ~hq ~0�q ~Oq ~(<q ~�q ~JSq ~��q ~d�q ~p q ~�q ~�q ~�q ~�$q ~�q ~6q ~3q ~Pq ~j.q ~(q ~[:q ~�q ~ttq ~ q ~#q ~ALq ~v�q ~x�q ~gq ~Imq ~�q ~$]q ~t�q ~/�q ~=<q ~Vq ~�q ~r�q ~�q ~�q ~N�q ~*jq ~l�q ~[�q ~r�q ~N$q ~?Dq ~?q ~!q ~*�q ~�q ~=�q ~T�q ~H�q ~O�q ~4�q ~`�q ~Uq ~yq ~GSq ~7;q ~3�q ~�q ~�q ~%�q ~%�q ~Pq ~-Zq ~dq ~$�q ~1q ~��q ~b>q ~#�q ~(uq ~c�q ~'q ~��q ~X�q ~,iq ~H�q ~Shq ~+�q ~�q ~(�q ~qq ~%]q ~R#q ~$q ~]uq ~9Lq ~q ~Bq ~t�q ~�q ~*]q ~��q ~��q ~Oq ~p�q ~�q ~3`q ~��q ~rq ~uQq ~b�q ~��q ~	�q ~9iq ~|�q ~�q ~s�q ~gq ~,�q ~k\q ~�q ~��q ~_q ~�q ~x�q ~9?q ~bq ~yq ~2pq ~�q ~�^q ~S�q ~`�q ~PRq ~�q ~�\q ~>�q ~��q ~V�q ~8q ~* q ~V�q ~@Cq ~
q ~Wmq ~G`q ~�q ~_q ~A�q ~E�q ~�Fq ~�q ~?�q ~q ~aq ~T�q ~/q ~>�q ~p�q ~L�q ~��q ~F<q ~I�q ~��q ~�q ~Iq ~��q ~\�q ~Z�q ~q ~@�q ~q ~g\q ~Gq ~�.q ~8�q ~:0q ~3mq ~CDq ~r�q ~�9q ~�q ~�$q ~�q ~��q ~f�q ~oRq ~"nq ~��q ~�Iq ~��q ~0�q ~BRq ~�q ~"�q ~��q ~Y�q ~Qgq ~�q ~w�q ~@&q ~jq ~:�q ~Z�q ~x<q ~1�q ~4�q ~.�q ~uq ~%q ~ hq ~]hq ~:Jq ~�q ~i1q ~�7q ~%�q ~��q ~[�q ~t�q ~�q ~<�q ~4�q ~8q ~X�q ~4$q ~��q ~n�q ~%yq ~O�q ~h�q ~Q=q ~��q ~4�q ~gq ~vq ~lfq ~�q ~q ~��q ~4�q ~AYq ~ yq ~$1q ~U�q ~Rsq ~u�q ~'�q ~M�q ~2�q ~�q ~�q ~#+q ~�q ~��q ~�q ~(�q ~�q ~u�q ~*q ~�q ~)@q ~0q ~=q ~�q ~�vq ~Rfq ~.q ~Yq ~�q ~5�q ~vq ~Q�q ~'�q ~�q ~C	q ~l*q ~mq ~��q ~dmq ~iSq ~Uq ~|�q ~�q ~)Mq ~zq ~Ehq ~[q ~
q ~v�q ~R�q ~`q ~KEq ~6q ~D�q ~-q ~�q ~g�q ~]Nq ~=�q ~?q ~w�q ~Aq ~W`q ~u{q ~/�q ~v�q ~zKq ~�&q ~@�q ~':q ~�q ~TIq ~F�q ~)"q ~<�q ~`�q ~~q ~	�q ~�q ~MIq ~��q ~�Oq ~�Mq ~��q ~pYq ~_�q ~?\q ~�q ~H2q ~	�q ~(/q ~�1q ~�Nq ~
�q ~*/q ~beq ~�gq ~6�q ~��q ~��q ~k�q ~��q ~[q ~"�q ~Fq ~Kq ~k�q ~jEq ~:dq ~vMq ~,�q ~X_q ~�q ~=q ~��q ~��q ~G/q ~�q ~|q ~<uq ~,q ~7�q ~>cq ~Mq ~S�q ~$�q ~aTq ~}�q ~1 q ~Yq ~;�q ~rq ~�Jq ~,@q ~#tq ~h�q ~&�q ~�q ~�q ~cq ~�q ~�q ~`iq ~YEq ~	@q ~Y�q ~N>q ~~�q ~g�q ~B�q ~_�q ~3�q ~A�q ~p/q ~#�q ~q ~�q ~��q ~�q ~zq ~Q�q ~K8q ~aq ~tgq ~1�q ~dSq ~&9q ~Gzq ~Xlq ~�~q ~m�q ~q ~a�q ~�q ~+�q ~?7q ~Nvq ~�]q ~��q ~Y+q ~;�q ~(�q ~Oxq ~ �q ~6�q ~7q ~��q ~]�q ~k5q ~J�q ~&q ~8wq ~f�q ~
Aq ~y�q ~ Tq ~[+q ~ffq ~RLq ~�sq ~I�q ~Qq ~oEq ~\Kq ~=Yq ~,�q ~n�q ~ZTq ~�q ~7�q ~}Yq ~B�q ~�Rq ~_�q ~;pq ~#q ~^�q ~qNq ~ �q ~aq ~��q ~�q ~fsq ~1}q ~I`q ~�q ~}�q ~wq ~~Aq ~0q ~emq ~�q ~[q ~"~q ~y^q ~�Qq ~Fq ~W�q ~E[q ~SAq ~xwq ~`�q ~q ~�*q ~jnq ~�q ~5q ~!q ~H�q ~�q ~��q ~/�q ~P�q ~$�q ~nq ~�q ~b�q ~H�q ~[�q ~t�q ~9�q ~b�q ~�q ~Uq ~�q ~�q ~�q ~��q ~q ~��q ~$�q ~�_q ~>Vq ~�{q ~&q ~�Dq ~>�q ~6�q ~r�q ~p�q ~}�q ~Myq ~~�q ~!�q ~y�q ~%q ~��q ~v�q ~�q ~Gq ~&�q ~�q ~-tq ~Uq ~]�q ~�q ~i�q ~�q ~f"q ~�q ~)rq ~7Lq ~�q ~-�q ~HLq ~)/q ~<�q ~P_q ~U�q ~9�q ~R2q ~~'q ~q�q ~lIq ~@�q ~28q ~�q ~oq ~�)q ~sAq ~#�q ~��q ~m1q ~ykq ~aaq ~6�q ~Eq ~H�q ~V�q ~Wq ~y�q ~n�q ~Yq ~fq ~(hq ~2q ~M(q ~�q ~9�q ~�2q ~	q ~zq ~]4q ~�q ~.q ~vwq ~lYq ~r7q ~y�q ~dFq ~.�q ~f�q ~~�q ~��q ~d�q ~>q ~q�q ~#�q ~q ~Oq ~m>q ~xq ~d�q ~K�q ~�q ~aGq ~��q ~q ~\q ~8q ~*�q ~}�q ~wxq ~M�q ~:=q ~ >q ~!Dq ~T�q ~Cq ~(Yq ~j�q ~t�q ~&�q ~u�q ~U�q ~]q ~Bq ~�q ~?�q ~hvq ~3Sq ~T�q ~+3q ~�q ~�q ~bvq ~^q ~��q ~&,q ~{�q ~~�q ~bKq ~kq ~Vwq ~&Fq ~Kiq ~�q ~gOq ~�q ~meq ~�q ~ �q ~4Mq ~6�q ~=q ~�@q ~�bq ~bXq ~M�q ~E�q ~�q ~%q ~=q ~<�q ~_�q ~m$q ~+`q ~	tq ~Xq ~_@q ~tZq ~FIq ~>q ~N�q ~/tq ~9%q ~4q ~i�q ~6gq ~$$q ~�8q ~F/q ~e�q ~l�q ~Ngq ~�q ~hXq ~s�q ~&�q ~Ueq ~xq ~�q ~C�q ~l:q ~\�q ~Eq ~T�q ~c�q ~#�q ~.Xq ~�q ~w�q ~�yq ~!Sq ~A�q ~P�q ~/�q ~a(q ~(�q ~+�q ~-Iq ~cq ~P+q ~��q ~�q ~K�q ~$�q ~P�q ~Gmq ~?�q ~G�q ~��q ~*�q ~8�q ~\�q ~ �q ~'�q ~C�q ~S�q ~t q ~W�q ~T�q ~�rq ~e�q ~6q ~<Vq ~Y_q ~Zq ~zgq ~"�q ~q�q ~ �q ~j�q ~qAq ~h�q ~/"q ~e�q ~kq ~y�q ~n�q ~Uq ~��q ~^<q ~A�q ~"�q ~3�q ~P�q ~7�q ~h�q ~y(q ~fq ~\5q ~<
q ~;�q ~!q ~|�q ~d�q ~|q ~$Pq ~A;q ~=nq ~6q ~s�q ~�q ~B�q ~��q ~+q ~d�q ~��q ~l�q ~_�q ~mXq ~�q ~q ~g�q ~�Rq ~-�q ~5�q ~�q ~,&q ~
�q ~��q ~�q ~s�q ~�~q ~,3q ~4gq ~z�q ~�q ~^�q ~VNq ~��q ~��q ~QWq ~2�q ~5�q ~�q ~G�q ~	q ~q ~�q ~; q ~K\q ~�Kq ~"8q ~|�q ~Sq ~d|q ~q ~��q ~�q ~�q ~J�q ~��q ~�Iq ~c�q ~�q ~}"q ~p�q ~=�q ~w�q ~jaq ~w�q ~W�q ~�q ~+q ~��q ~/�q ~v]q ~�q ~q ~<eq ~1�q ~#q ~x�q ~"�q ~�q ~SNq ~!#q ~Nq ~m�q ~��q ~Mjq ~iq ~W'q ~j�q ~��q ~Mq ~y5q ~@6q ~7!q ~g(q ~{�q ~@q ~1q ~.Gq ~r�q ~.eq ~	Qq ~0@q ~(q ~��q ~#q ~��q ~Qtq ~b�q ~l�q ~rrq ~N�q ~U�q ~%�q ~}q ~B�q ~o+q ~F�q ~*�q ~?�q ~(�q ~3�q ~;Gq ~�q ~//q ~)q ~0zq ~L�q ~4Zq ~>�q ~�q ~�q ~jq ~"�q ~�q ~Hq ~tq ~Wq ~{�q ~%?q ~��q ~��q ~/q ~<�q ~��q ~�q ~/q ~Urq ~ �q ~lq ~B"q ~4�q ~?�q ~?�q ~cVq ~~�q ~�q ~�q ~]�q ~?lq ~(q ~ �q ~q ~H�q ~��q ~V]q ~Qq ~c�q ~xq ~;�q ~A�q ~�q ~]�q ~ �q ~XRq ~Z�q ~�xq ~C�q ~�q ~u�q ~aq ~:�q ~K�q ~s�q ~cq ~8q ~U;q ~)eq ~8jq ~��q ~|!q ~v�q ~rq ~&�q ~Fq ~S'q ~6q ~'�q ~rq ~d/q ~�q ~6q ~U�q ~_~q ~H�q ~%q ~S[q ~X�q ~Biq ~J�q ~�/q ~O	q ~\�q ~��q ~v�q ~ �q ~Rq ~'�q ~m�q ~Kyq ~e�q ~*{q ~��q ~BEq ~z�q ~_�q ~q ~�q ~n�q ~+mq ~g�q ~�q ~q ~Oiq ~�q ~�q ~T�q ~{�q ~u*q ~Q�q ~�q ~�q ~Mq ~[�q ~Jq ~<Gq ~Fq ~z�q ~h.q ~ �q ~t>q ~2Vq ~6Jq ~!�q ~��q ~Lfq ~��q ~&dq ~v�q ~�q ~Zq ~ipq ~v@q ~$q ~eOq ~5�q ~H�q ~MZq ~7Yq ~>q ~C�q ~A�q ~Zaq ~W�q ~Fq ~G�q ~q ~%�q ~kq ~� q ~{~q ~j�q ~�q ~!�q ~`(q ~hq ~gq ~$�q ~8(q ~��q ~z$q ~bq ~,�q ~kvq ~S�q ~Q�q ~[rq ~�q ~%q ~N�q ~�q ~��q ~88q ~)�q ~��q ~�q ~H�q ~M�q ~�q ~\q ~"(q ~sQq ~@{q ~O2q ~�q ~�q ~Eq ~~q ~xjq ~�q ~�q ~-�q ~mq ~;'q ~{dq ~�q ~1�q ~7�q ~�q ~Gq ~Jxq ~q ~Tq ~�vq ~Yq ~"q ~<q ~&�q ~��q ~�q ~+�q ~0`q ~[Gq ~�q ~`\q ~�_q ~r�q ~3Fq ~@q ~>q ~�q ~��q ~N�q ~_q ~U�q ~��q ~Dq ~m�q ~wQq ~= q ~�q ~o�q ~\�q ~,�q ~p�q ~�q ~~�q ~D�q ~!`q ~l�q ~��q ~R�q ~�Wq ~��q ~�q ~>�q ~4q ~�q ~2�q ~]�q ~aq ~�q ~wDq ~`�q ~�_q ~.+q ~NMq ~I�q ~13q ~ q ~�?q ~H�q ~~�q ~C&q ~0Pq ~�;q ~^�q ~��q ~q ~
Sq ~F�q ~v0q ~�q ~�fq ~0�q ~kq ~��q ~M�q ~'�q ~N�q ~��q ~�q ~h�q ~�q ~��q ~[eq ~�q ~X�q ~�q ~��q ~/q ~�q ~=�q ~OOq ~o�q ~~q ~_dq ~k�q ~2'q ~/�q ~f/q ~�q ~sq ~gBq ~�6q ~?�q ~pfq ~�q ~�"q ~Eq ~'*q ~g�q ~CQq ~<�q ~�q ~q ~quq ~]Aq ~J�q ~fIq ~�q ~'�q ~n&q ~j�q ~Aq ~vq ~
�q ~G<q ~=�q ~�q ~q ~iq ~P�q ~o�q ~d�q ~�cq ~wq ~Trq ~ �q ~�dq ~Y�q ~yq ~U�q ~:�q ~
�q ~vq ~a�q ~�#q ~{'q ~|�q ~E�q ~z�q ~�q ~w�q ~��q ~{�q ~V"q ~X�q ~Z�q ~�q ~cIq ~aq ~�q ~<�q ~O#q ~O@q ~S}q ~8�q ~n�q ~X�q ~^Kq ~�q ~y�q ~�q ~�q ~��q ~X�q ~{�q ~`�q ~1�q ~M8q ~4q ~m�q ~�q ~q ~,q ~:~q ~�q ~}nq ~\q ~ /q ~Kq ~�q ~a�q ~"q ~%/q ~�q ~e�q ~�Zq ~K�q ~	�q ~�q ~@Pq ~��q ~+�q ~U�q ~�q ~N�q ~|.q ~C3q ~y�q ~(q ~:�q ~K�q ~[q ~:�q ~L�q ~x"q ~Jq ~b�q ~�q ~&�q ~8�q ~4q ~Hwq ~|[q ~9q ~~hq ~#Iq ~|=q ~Q�q ~-q ~D-q ~_Oq ~	
q ~6Zq ~��q ~��q ~][q ~PEq ~c�q ~@�q ~`q ~%"q ~��q ~*Kq ~nNq ~�^q ~�q ~RYq ~&q ~I�q ~Zq ~~�q ~��q ~b�q ~;6q ~F�q ~c�q ~mrq ~T�q ~p�q ~j�q ~v�q ~gq ~C�q ~U�q ~��q ~R�q ~Vq ~B�q ~;�q ~t1q ~s^q ~W�q ~/Zq ~vq ~ +q ~z�q ~h�q ~W4q ~r�q ~TXq ~G�q ~Cq ~�q ~
tq ~WAq ~Gq ~>q ~f�q ~L2q ~#q ~�q ~z�q ~!�q ~�q ~)�q ~�q ~?*q ~)�q ~��q ~�q ~]'q ~�q ~C�q ~'q ~
0q ~Tq ~39q ~�q ~1Dq ~<1q ~0�q ~J�q ~�uq ~mq ~}�q ~Q�q ~_�q ~��q ~��q ~x�q ~�q ~pq ~�~q ~��q ~Oq ~E�q ~*�q ~Tq ~rq ~3�q ~�q ~uq ~�q ~�q ~�=q ~yQq ~{q ~
cq ~
q ~Lq ~y�q ~|�q ~�q ~{Jq ~ooq ~pq ~'\q ~3q ~D�q ~nzq ~5�q ~yDq ~5�q ~o�q ~vq ~��q ~Mq ~{qq ~�rq ~Hq ~>�q ~"�q ~.:q ~qq ~��q ~eq ~eq ~m�q ~GFq ~R�q ~E�q ~ICq ~v�q ~q ~q ~4�q ~l�q ~_�q ~�q ~~[q ~%�q ~M�q ~�q ~e>q ~�q ~9�q ~�q ~
�q ~B8q ~+q ~)�q ~K)q ~�q ~5Dq ~2q ~\�q ~��q ~�q ~�)q ~R?q ~zwq ~�q ~D�q ~_3q ~`�q ~�;q ~4�q ~s�q ~�q ~`Bq ~e�q ~iFq ~<�q ~8q ~��q ~%�q ~L�q ~?yq ~wq ~�fq ~5q ~c�q ~6�q ~xKq ~Zq ~e�q ~)�q ~c/q ~�q ~.�q ~<�q ~�q ~Gq ~kOq ~�q ~��q ~�\q ~Q#q ~2q ~G�q ~��q ~^�q ~Frq ~Byq ~x�q ~Asq ~+&q ~w�q ~9q ~T�q ~�3q ~'q ~k�q ~(�q ~e�q ~q ~z�q ~`Oq ~Q0q ~�q ~z�q ~q ~rTq ~@q ~�q ~[�q ~4�q ~%Lq ~>q ~g5q ~R�q ~~q ~�7q ~�q ~}/q ~g�q ~��q ~>&q ~xq ~q ~]q ~|q ~Fcq ~ "q ~zq ~sq ~jRq ~�q ~/gq ~\[q ~0/q ~�qq ~ezq ~S q ~��q ~�[q ~b�q ~q�q ~�q ~�q ~#�q ~;cq ~�q ~rDq ~��q ~]�q ~psq ~c�q ~��q ~G�q ~\�q ~^�q ~a�q ~)�q ~�Qq ~l�q ~�"q ~�q ~L�q ~�q ~hKq ~�q ~{q ~1aq ~j!q ~H?q ~h�q ~:#q ~g�q ~Mq ~1�q ~A�q ~��q ~.�q ~i�q ~S4q ~.�q ~q[q ~i�q ~{�q ~7�q ~/�q ~w(q ~4tq ~=�q ~:q ~7q ~E�q ~hq ~%�q ~�lq ~9�q ~�>q ~Jq ~��q ~Nq ~7�q ~��q ~�Yq ~%jq ~q ~Jq ~m�q ~@�q ~��q ~^sq ~E3q ~:qq ~8q ~[�q ~Xq ~x�q ~�Xq ~Lsq ~:�q ~	�q ~Uq ~h�q ~zq ~�q ~9zq ~�q ~^�q ~�qq ~*<q ~;�q ~Nq ~�jq ~�,q ~+q ~lwq ~ �q ~W q ~U.q ~�q ~i�q ~��q ~Xq ~-�q ~lq ~��q ~w�q ~I)q ~�q ~#Vq ~Gq ~�q ~uq ~.�q ~b"q ~�q ~S�q ~5)q ~C�q ~�kq ~r�q ~lq ~ctq ~�q ~`5q ~j}q ~cq ~}{q ~��q ~o�q ~'mq ~ q ~wkq ~Z�q ~q ~D�q ~q ~Y�q ~5�q ~	�q ~.�q ~W�q ~FVq ~vjq ~!q ~,�q ~�q ~5^q ~6�q ~^�q ~Z�q ~�Yq ~qq ~Tq ~S�q ~b�q ~g�q ~��q ~+@q ~&tq ~B�q ~�q ~e"q ~-�q ~i$q ~0q ~�3q ~Pq ~��q ~V?q ~h;q ~w7q ~q ~0�q ~�Wq ~Z�q ~u7q ~_q ~ lq ~,Oq ~Hq ~}<q ~�tq ~P�q ~w�q ~|hq ~R�q ~q ~
�q ~i�q ~��q ~�Eq ~Y�q ~�q ~*�q ~L�q ~Wzq ~q�q ~qq ~Oq ~�lq ~?�q ~6q ~,\q ~J�q ~ �q ~E#q ~kiq ~[�q ~��q ~a�q ~�q ~*�q ~�q ~Sq ~j�q ~g�q ~�yq ~q ~�q ~a8q ~�,q ~W�q ~�q ~y�q ~Kq ~�q ~�hq ~F�q ~�q ~^q ~k�q ~8�q ~#cq ~+�q ~V1q ~'q ~	1q ~H%q ~��q ~-9q ~W�q ~S�q ~u�q ~7�q ~s�q ~eq ~�
q ~	�q ~N�q ~f�q ~|Jq ~��q ~��q ~G�q ~ Oq ~a�q ~B�q ~D�q ~Z�q ~=�q ~5�q ~I�q ~x/q ~cq ~�q ~gq ~�q ~t�q ~�q ~6=q ~<�q ~hq ~)�q ~Wq ~Iq ~�q ~Jbq ~)�q ~�q ~�q ~��q ~Bq ~@�q ~=q ~�#q ~,q ~m�q ~{�q ~Nq ~3�q ~<q ~'�q ~�!q ~"Hq ~0mq ~}�q ~�q ~.�q ~ |q ~-�q ~o_q ~f�q ~R�q ~��q ~@_q ~]�q ~Afq ~mq ~�q ~J�q ~?q ~&Sq ~I~q ~,�q ~!�q ~q ~�Rq ~Eq ~`
q ~q'q ~'~q ~}Iq ~|q ~Pq ~=Iq ~7�q ~�q ~�q ~o�q ~�
q ~D<q ~u�q ~�*q ~I6q ~,vq ~��q ~�Jq ~�"q ~gq ~d`q ~dq ~n�q ~3�q ~L%q ~ q ~zZq ~4q ~h!q ~ _q ~�
q ~pq ~�q ~Dq ~�@q ~)q ~q ~apq ~
�q ~1Tq ~NZq ~i`q ~-gq ~/�q ~P�q ~|�q ~@�q ~Wq ~*q ~`�q ~J9q ~^/q ~�$q ~J,q ~�iq ~2�q ~��q ~aq ~V�q ~t�q ~Teq ~tq ~oq ~|q ~<$q ~P8q ~Z�q ~L�q ~f<q ~L?q ~X�q ~zq ~~uq ~'Kq ~unq ~\�q ~XEq ~"
q ~JFq ~�q ~��q ~z1q ~UJq ~�q ~4�q ~K�q ~��q ~O�q ~>7q ~C^q ~^�q ~uaq ~�q ~YRq ~	q ~Cxq ~�q ~��q ~��q ~\hq ~N1q ~}�q ~D^q ~��q ~a�q ~7�q ~s�q ~ZDq ~Y�q ~gvq ~oq ~C�q ~|�q ~:�q ~�Fq ~�q ~O�q ~�q ~9�q ~�q ~8�q ~Y�q ~V�q ~
�q ~?�q ~w^q ~�q ~(Iq ~�q ~w�q ~\�q ~iq ~{4q ~dq ~:q ~0�q ~>Gq ~yxq ~V�q ~#�q ~$q ~*q ~iq ~#;q ~p<q ~�q ~QJq ~��q ~A.q ~��q ~D�xq ~��sq ~��w   ?@     q ~�{xq ~=ksq ~��w   ?@     q ~Iq ~j;q ~B_q ~"aq ~=fq ~ �xq ~[�sq ~��w   ?@     q ~[�xq ~_asq ~��w   ?@     q ~��q ~��q ~_\q ~v�q ~h�q ~�*q ~q ~R
q ~q ~�Hq ~Mxq ~P�sq ~��w   ?@     q ~P�q ~d<xq ~Asq ~��w   @?@     -q ~e�q ~~Nq ~n_q ~��q ~�/q ~b�q ~qq ~R�q ~��q ~`�q ~V�q ~�q ~?Qq ~b�q ~q ~iq ~,�q ~oq ~2q ~p�q ~$Bq ~o q ~Z,q ~�q ~sxq ~5�q ~heq ~1q ~eq ~>�q ~%�q ~+q ~;q ~�q ~$�q ~h�q ~q ~qq ~��q ~KRq ~�q ~WNq ~Aq ~o8q ~��xq ~	)sq ~��w   ?@     
q ~	q ~�q ~5{q ~O�q ~t�q ~�q ~��q ~u�q ~Doq ~Vjxq ~n�sq ~��w   @?@     q ~Euq ~Yq ~M�q ~1�q ~�q ~7q ~�<q ~U�q ~�q ~Pyq ~(�q ~Q�q ~�kq ~.�q ~n�q ~��q ~��q ~I�q ~�sq ~�q ~-�q ~�Sq ~9 q ~5q ~}�q ~Q�q ~xxq ~�sq ~��w    ?@     q ~W�q ~��q ~}fq ~@q ~�q ~S�q ~M�q ~]q ~i>q ~-q ~E�q ~�q ~}�q ~p�q ~Aq ~��q ~56xq ~`"sq ~��w   ?@     q ~`xq ~m�sq ~��w   ?@     q ~mxq ~�'sq ~��w   ?@     q ~jq ~>yq ~�.q ~�q ~�"xq ~t.sq ~��w   ?@     q ~t)q ~i�xq ~Nsq ~��w   ?@     q ~<q ~&�q ~�xxsq ~ C?@     w       q ~��sq ~��w   ?@     q ~��q ~��xq ~�9sq ~��w   ?@     	q ~��q ~��q ~��q ~��q ~��q ~�4q ~��q ~�!q ~�nxq ~�6sq ~��w   ?@     q ~�1xq ~�!sq ~��w    ?@     q ~��q ~�Iq ~�iq ~�Sq ~�q ~�q ~��q ~��q ~�q ~��q ~��q ~��q ~��q ~��q ~��q ~�q ~�q ~�qq ~�Gq ~�q ~�xq ~�dsq ~��w   ?@     q ~�dq ~�3q ~�_xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��q ~��xq ~�Ksq ~��w   ?@     q ~�Fxq ~�:sq ~��w   ?@     q ~�5q ~��q ~�xq ~��sq ~��w   ?@     q ~��xq ~�Osq ~��w   ?@     	q ~��q ~��q ~�q ~��q ~�Yq ~��q ~�Jq ~�q ~��xq ~�$sq ~��w   ?@     	q ~��q ~�0q ~��q ~�Dq ~�8q ~�rq ~�aq ~�q ~�+xq ~��sq ~��w   ?@     q ~��q ~��q ~��xq ~�Zsq ~��w   ?@     q ~��q ~�{q ~��q ~�Uq ~�Wq ~�6q ~��q ~��q ~�Vq ~��q ~��xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~��xq ~��sq ~��w   ?@     q ~�8q ~��q ~�q ~��xq ~�rsq ~��w   ?@     q ~�mq ~��xq ~�sq ~��w   ?@     q ~�xxsr 9edu.cornell.cs.nlp.spf.base.hashvector.FastTreeHashVector;��tQ57� L valuest 0Lit/unimi/dsi/fastutil/objects/Object2DoubleMap;xpsr 5it.unimi.dsi.fastutil.objects.Object2DoubleAVLTreeMap�7y�J| I countL storedComparatort Ljava/util/Comparator;xr <it.unimi.dsi.fastutil.objects.AbstractObject2DoubleSortedMap�c����  xr 6it.unimi.dsi.fastutil.objects.AbstractObject2DoubleMap�o��K<z  xr ;it.unimi.dsi.fastutil.objects.AbstractObject2DoubleFunction�o��K<z D defRetValuexp          �psq ~��WD�t DYNSKIPppppw��      sq ~��W�"�q ~ t LEXt 0t 0pw        sq ~��W���q ~ q ~�9t 0t 18pw@5oz�G�sq ~��W�#4q ~ q ~�9t 0t 3pw        sq ~��W�#�q ~ q ~�9t 0t 6pw        sq ~��W�&�q ~ q ~�9t 1t 1pw@$      sq ~��W�!q ~ q ~�9t 10t 11pw@$      sq ~��W�%Sq ~ q ~�9t 10t 25pw@%���}B�sq ~��W�0�q ~ q ~�9t 10t 57pw        sq ~��Zw0�q ~ q ~�9t 100t 27pw@-�|���sq ~��Zw?q ~ q ~�9t 100t 60pw@$�1��$sq ~�ή�q ~ q ~�9t 1000t 61pw        sq ~�ή��q ~ q ~�9t 1000t 84pw@F�U�i�sq ~�ή��q ~ q ~�9t 1001t 61pw        sq ~�ή��q ~ q ~�9t 1001t 84pw@5oz�G�sq ~�ή�|q ~ q ~�9t 1002t 84pw@5oz�G�sq ~�ή�^q ~ q ~�9t 1003t 61pw        sq ~�ή�=q ~ q ~�9t 1003t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1004t 84pw@@�鹙�sq ~�ή�q ~ q ~�9t 1005t 75pw        sq ~�ή��q ~ q ~�9t 1005t 84pw@$      sq ~�ή��q ~ q ~�9t 1006t 84pw@@�鹙�sq ~�ή�bq ~ q ~�9t 1007t 61pw        sq ~�ή�Aq ~ q ~�9t 1007t 84pw@@�鹙�sq ~�ή�`q ~ q ~�9t 1008t 75pw        sq ~�ή�q ~ q ~�9t 1008t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1009t 61pw        sq ~�ή��q ~ q ~�9t 1009t 84pw@@�鹙�sq ~��ZwG�q ~ q ~�9t 101t 79pw@@�鹙�sq ~�ήYq ~ q ~�9t 1010t 84pw@5oz�G�sq ~�ήxq ~ q ~�9t 1011t 75pw        sq ~�ήq ~ q ~�9t 1011t 84pw@5oz�G�sq ~�ή!�q ~ q ~�9t 1012t 84pw@5oz�G�sq ~�ή%�q ~ q ~�9t 1013t 84pw@F�U�i�sq ~�ή!~q ~ q ~�9t 1014t 61pw        sq ~�ή)]q ~ q ~�9t 1014t 84pw@F�U�i�sq ~�ή-q ~ q ~�9t 1015t 84pw@$      sq ~�ή0�q ~ q ~�9t 1016t 84pw@5oz�G�sq ~�ή4�q ~ q ~�9t 1017t 84pw@5oz�G�sq ~�ή4�q ~ q ~�9t 1018t 75pw        sq ~�ή8aq ~ q ~�9t 1018t 84pw@5oz�G�sq ~�ή4Cq ~ q ~�9t 1019t 61pw        sq ~�ή<"q ~ q ~�9t 1019t 84pw@$      sq ~��ZwNq ~ q ~�9t 102t 80pw@5oz�G�sq ~��ZwNoq ~ q ~�9t 102t 83pw@5oz�G�sq ~�ή��q ~ q ~�9t 1020t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1021t 75pw        sq ~�ή�yq ~ q ~�9t 1021t 84pw@5oz�G�sq ~�ή�[q ~ q ~�9t 1022t 61pw        sq ~�ή�:q ~ q ~�9t 1022t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1023t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1024t 84pw@$      sq ~�ή�}q ~ q ~�9t 1025t 84pw@$      sq ~�ή�_q ~ q ~�9t 1026t 61pw        sq ~�ή�>q ~ q ~�9t 1026t 84pw@$      sq ~�ή�]q ~ q ~�9t 1027t 75pw        sq ~�ή��q ~ q ~�9t 1027t 84pw@$      sq ~�ή��q ~ q ~�9t 1028t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1029t 61pw        sq ~�ή��q ~ q ~�9t 1029t 84pw@$      sq ~��ZwQ�q ~ q ~�9t 103t 81pw@@�鹙�sq ~�ήq ~ q ~�9t 1030t 84pw@F�U�i�sq ~�ή��q ~ q ~�9t 1031t 61pw        sq ~�ή�q ~ q ~�9t 1031t 84pw@$      sq ~�ή
�q ~ q ~�9t 1032t 84pw@5oz�G�sq ~�ή{q ~ q ~�9t 1033t 61pw        sq ~�ήZq ~ q ~�9t 1033t 84pw@5oz�G�sq ~�ήq ~ q ~�9t 1034t 84pw@@�鹙�sq ~�ή�q ~ q ~�9t 1035t 61pw        sq ~�ή�q ~ q ~�9t 1035t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1036t 61pw        sq ~�ή�q ~ q ~�9t 1036t 84pw@5oz�G�sq ~�ή^q ~ q ~�9t 1037t 84pw@5oz�G�sq ~�ή!q ~ q ~�9t 1038t 84pw@$      sq ~�ήq ~ q ~�9t 1039t 61pw        sq ~�ή$�q ~ q ~�9t 1039t 84pw@F�U�i�sq ~��ZwU�q ~ q ~�9t 104t 82pw@$      sq ~�ήo�q ~ q ~�9t 1040t 61pw        sq ~�ήwvq ~ q ~�9t 1040t 84pw@$      sq ~�ή{7q ~ q ~�9t 1041t 84pw@5oz�G�sq ~�ήwq ~ q ~�9t 1042t 61pw        sq ~�ή~�q ~ q ~�9t 1042t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1043t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1044t 75pw        sq ~�ή�zq ~ q ~�9t 1044t 84pw@F�U�i�sq ~�ή�\q ~ q ~�9t 1045t 61pw        sq ~�ή�;q ~ q ~�9t 1045t 84pw@$      sq ~�ή�q ~ q ~�9t 1046t 61pw        sq ~�ή��q ~ q ~�9t 1046t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1047t 75pw        sq ~�ή��q ~ q ~�9t 1047t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1048t 75pw        sq ~�ή�~q ~ q ~�9t 1048t 84pw@@�鹙�sq ~�ή�?q ~ q ~�9t 1049t 84pw@$      sq ~��ZwY�q ~ q ~�9t 105t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1050t 84pw@@�鹙�sq ~�ή�q ~ q ~�9t 1051t 84pw@5oz�G�sq ~�ή�xq ~ q ~�9t 1052t 61pw        sq ~�ή�Wq ~ q ~�9t 1052t 84pw@F�U�i�sq ~�ή�vq ~ q ~�9t 1053t 75pw        sq ~�ή�q ~ q ~�9t 1053t 84pw@5oz�G�sq ~�ή�7q ~ q ~�9t 1054t 75pw        sq ~�ή��q ~ q ~�9t 1054t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1055t 61pw        sq ~�ή��q ~ q ~�9t 1055t 84pw@$      sq ~�ή�|q ~ q ~�9t 1056t 61pw        sq ~�ή	[q ~ q ~�9t 1056t 84pw@5oz�G�sq ~�ή�=q ~ q ~�9t 1057t 61pw        sq ~�ή	q ~ q ~�9t 1057t 84pw@5oz�G�sq ~�ή	;q ~ q ~�9t 1058t 75pw        sq ~�ή		�q ~ q ~�9t 1058t 84pw@$      sq ~�ή	�q ~ q ~�9t 1059t 61pw        sq ~�ή	�q ~ q ~�9t 1059t 84pw@$      sq ~��Zw]�q ~ q ~�9t 106t 84pw@$      sq ~�ή	\�q ~ q ~�9t 1060t 75pw        sq ~�ή	`4q ~ q ~�9t 1060t 84pw@F�U�i�sq ~�ή	\q ~ q ~�9t 1061t 61pw        sq ~�ή	c�q ~ q ~�9t 1061t 84pw@F�U�i�sq ~�ή	dq ~ q ~�9t 1062t 75pw        sq ~�ή	g�q ~ q ~�9t 1062t 84pw@5oz�G�sq ~�ή	c�q ~ q ~�9t 1063t 61pw        sq ~�ή	kwq ~ q ~�9t 1063t 84pw@5oz�G�sq ~�ή	gYq ~ q ~�9t 1064t 61pw        sq ~�ή	o8q ~ q ~�9t 1064t 84pw@F�U�i�sq ~�ή	kq ~ q ~�9t 1065t 61pw        sq ~�ή	r�q ~ q ~�9t 1065t 84pw@@�鹙�sq ~�ή	n�q ~ q ~�9t 1066t 61pw        sq ~�ή	v�q ~ q ~�9t 1066t 84pw@@�鹙�sq ~�ή	r�q ~ q ~�9t 1067t 61pw        sq ~�ή	z{q ~ q ~�9t 1067t 84pw@#�K`�Esq ~�ή	~<q ~ q ~�9t 1068t 84pw@$      sq ~�ή	~[q ~ q ~�9t 1069t 75pw        sq ~�ή	��q ~ q ~�9t 1069t 84pw@F�U�i�sq ~��ZwYtq ~ q ~�9t 107t 61pw        sq ~��ZwaSq ~ q ~�9t 107t 84pw@@�鹙�sq ~�ή	��q ~ q ~�9t 1070t 75pw        sq ~�ή	ԓq ~ q ~�9t 1070t 84pw@@�鹙�sq ~�ή	Բq ~ q ~�9t 1071t 75pw        sq ~�ή	�Tq ~ q ~�9t 1071t 84pw@5oz�G�sq ~�ή	�6q ~ q ~�9t 1072t 61pw        sq ~�ή	�q ~ q ~�9t 1072t 84pw@@�鹙�sq ~�ή	��q ~ q ~�9t 1073t 61pw        sq ~�ή	��q ~ q ~�9t 1073t 84pw@5oz�G�sq ~�ή	�q ~ q ~�9t 1074t 84pw@@�鹙�sq ~�ή	�yq ~ q ~�9t 1075t 61pw        sq ~�ή	�Xq ~ q ~�9t 1075t 84pw@F�U�i�sq ~�ή	�q ~ q ~�9t 1076t 84pw@$      sq ~�ή	��q ~ q ~�9t 1077t 61pw        sq ~�ή	��q ~ q ~�9t 1077t 84pw@F�U�i�sq ~�ή	�q ~ q ~�9t 1078t 84pw@5oz�G�sq ~�ή	�\q ~ q ~�9t 1079t 84pw@$      sq ~��Zweq ~ q ~�9t 108t 84pw@@�鹙�sq ~�ή
EPq ~ q ~�9t 1080t 75pw        sq ~�ή
H�q ~ q ~�9t 1080t 84pw@5oz�G�sq ~�ή
Iq ~ q ~�9t 1081t 75pw        sq ~�ή
L�q ~ q ~�9t 1081t 84pw@@�鹙�sq ~�ή
L�q ~ q ~�9t 1082t 75pw        sq ~�ή
Ptq ~ q ~�9t 1082t 84pw@5oz�G�sq ~�ή
T5q ~ q ~�9t 1083t 84pw@@�鹙�sq ~�ή
TTq ~ q ~�9t 1084t 75pw        sq ~�ή
W�q ~ q ~�9t 1084t 84pw@5oz�G�sq ~�ή
[�q ~ q ~�9t 1085t 84pw@5oz�G�sq ~�ή
_xq ~ q ~�9t 1086t 84pw@@�鹙�sq ~�ή
[Zq ~ q ~�9t 1087t 61pw        sq ~�ή
c9q ~ q ~�9t 1087t 84pw@$      sq ~�ή
f�q ~ q ~�9t 1088t 84pw@$      sq ~�ή
j�q ~ q ~�9t 1089t 84pw@5oz�G�sq ~��Zwh�q ~ q ~�9t 109t 84pw@@�鹙�sq ~�ή
�Qq ~ q ~�9t 1090t 84pw@5oz�G�sq ~�ή
�q ~ q ~�9t 1091t 84pw@@�鹙�sq ~�ή
�1q ~ q ~�9t 1092t 75pw        sq ~�ή
��q ~ q ~�9t 1092t 84pw@$      sq ~�ή
��q ~ q ~�9t 1093t 61pw        sq ~�ή
Ȕq ~ q ~�9t 1093t 84pw@$      sq ~�ή
ȳq ~ q ~�9t 1094t 75pw        sq ~�ή
�Uq ~ q ~�9t 1094t 84pw@@�鹙�sq ~�ή
�q ~ q ~�9t 1095t 84pw@$      sq ~�ή
��q ~ q ~�9t 1096t 61pw        sq ~�ή
��q ~ q ~�9t 1096t 84pw@$      sq ~�ή
טq ~ q ~�9t 1097t 84pw@@�鹙�sq ~�ή
׷q ~ q ~�9t 1098t 75pw        sq ~�ή
�Yq ~ q ~�9t 1098t 84pw@5oz�G�sq ~�ή
�;q ~ q ~�9t 1099t 61pw        sq ~�ή
�q ~ q ~�9t 1099t 84pw@@�鹙�sq ~��W�$�q ~ q ~�9t 11t 12pw?�K�sq ~��W�%rq ~ q ~�9t 11t 16pw@$㼁���sq ~��W�(�q ~ q ~�9t 11t 23pw@-���%��sq ~��W�)qq ~ q ~�9t 11t 28pw��UQޥsq ~��W�)�q ~ q ~�9t 11t 29pw        sq ~��W�,xq ~ q ~�9t 11t 32pw�T<����Hsq ~��W�-Qq ~ q ~�9t 11t 39pw        sq ~��W�3�q ~ q ~�9t 11t 51pw        sq ~��Zw��q ~ q ~�9t 110t 75pw        sq ~��Zw�kq ~ q ~�9t 110t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1100t 61pw        sq ~�ή�{q ~ q ~�9t 1100t 84pw@$      sq ~�ή�<q ~ q ~�9t 1101t 84pw@$      sq ~�ή��q ~ q ~�9t 1102t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1103t 61pw        sq ~�ήȾq ~ q ~�9t 1103t 84pw@F�U�i�sq ~�ή�q ~ q ~�9t 1104t 84pw@5oz�G�sq ~�ή̞q ~ q ~�9t 1105t 75pw        sq ~�ή�@q ~ q ~�9t 1105t 84pw@#�ϗ�X�sq ~�ή�"q ~ q ~�9t 1106t 61pw        sq ~�ή�q ~ q ~�9t 1106t 84pw@F�U�i�sq ~�ή��q ~ q ~�9t 1107t 61pw        sq ~�ή��q ~ q ~�9t 1107t 84pw@@�鹙�sq ~�ήӤq ~ q ~�9t 1108t 61pw        sq ~�ήۃq ~ q ~�9t 1108t 84pw@$      sq ~�ή�eq ~ q ~�9t 1109t 61pw        sq ~�ή�Dq ~ q ~�9t 1109t 84pw@5oz�G�sq ~��Zw��q ~ q ~�9t 111t 75pw        sq ~��Zw�,q ~ q ~�9t 111t 84pw@F�U�i�sq ~�ή.8q ~ q ~�9t 1110t 75pw        sq ~�ή1�q ~ q ~�9t 1110t 84pw@$      sq ~�ή-�q ~ q ~�9t 1111t 61pw        sq ~�ή5�q ~ q ~�9t 1111t 84pw@$      sq ~�ή9\q ~ q ~�9t 1112t 84pw@5oz�G�sq ~�ή9{q ~ q ~�9t 1113t 75pw        sq ~�ή=q ~ q ~�9t 1113t 84pw@$      sq ~�ή8�q ~ q ~�9t 1114t 61pw        sq ~�ή@�q ~ q ~�9t 1114t 84pw@5oz�G�sq ~�ή@�q ~ q ~�9t 1115t 75pw        sq ~�ήD�q ~ q ~�9t 1115t 84pw@F�U�i�sq ~�ή@�q ~ q ~�9t 1116t 61pw        sq ~�ήH`q ~ q ~�9t 1116t 84pw@#��W�6sq ~�ήDBq ~ q ~�9t 1117t 61pw        sq ~�ήL!q ~ q ~�9t 1117t 84pw@F�U�i�sq ~�ήHq ~ q ~�9t 1118t 61pw        sq ~�ήO�q ~ q ~�9t 1118t 84pw@5oz�G�sq ~�ήK�q ~ q ~�9t 1119t 61pw        sq ~�ήS�q ~ q ~�9t 1119t 84pw@5oz�G�sq ~��Zw��q ~ q ~�9t 112t 84pw@$      sq ~�ή��q ~ q ~�9t 1120t 75pw        sq ~�ή�9q ~ q ~�9t 1120t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1121t 84pw@$      sq ~�ή�q ~ q ~�9t 1122t 75pw        sq ~�ή��q ~ q ~�9t 1122t 84pw@M]��%��sq ~�ή��q ~ q ~�9t 1123t 61pw����F�sq ~�ή�|q ~ q ~�9t 1123t 84pw@*j��0��sq ~�ή�=q ~ q ~�9t 1124t 84pw@F�U�i�sq ~�ή�\q ~ q ~�9t 1125t 75pw        sq ~�ή��q ~ q ~�9t 1125t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1126t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1127t 61pw        sq ~�ή��q ~ q ~�9t 1127t 84pw@5oz�G�sq ~�ή�Aq ~ q ~�9t 1128t 84pw@5oz�G�sq ~�ή�`q ~ q ~�9t 1129t 75pw        sq ~�ή�q ~ q ~�9t 1129t 84pw@5oz�G�sq ~��Zw�q ~ q ~�9t 113t 75pw        sq ~��ZwƮq ~ q ~�9t 113t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1130t 84pw@$��G74sq ~�ήzq ~ q ~�9t 1131t 61pw        sq ~�ήYq ~ q ~�9t 1131t 84pw@%�����ksq ~�ή"q ~ q ~�9t 1132t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1133t 61pw        sq ~�ή%�q ~ q ~�9t 1133t 84pw@5oz�G�sq ~�ή!�q ~ q ~�9t 1134t 61pw        sq ~�ή)�q ~ q ~�9t 1134t 84pw@@�鹙�sq ~�ή-]q ~ q ~�9t 1135t 84pw@@�鹙�sq ~�ή)?q ~ q ~�9t 1136t 61pw        sq ~�ή1q ~ q ~�9t 1136t 84pw@5oz�G�sq ~�ή4�q ~ q ~�9t 1137t 84pw@$      sq ~�ή8�q ~ q ~�9t 1138t 84pw@$      sq ~�ή4�q ~ q ~�9t 1139t 61pw        sq ~�ή<aq ~ q ~�9t 1139t 84pw@5oz�G�sq ~��Zwq ~ q ~�9t 114t 61pw        sq ~��Zw�oq ~ q ~�9t 114t 84pw@A96�XZsq ~�ή�Uq ~ q ~�9t 1140t 75pw        sq ~�ή��q ~ q ~�9t 1140t 84pw@@�鹙�sq ~�ή�q ~ q ~�9t 1141t 75pw        sq ~�ή��q ~ q ~�9t 1141t 84pw@$      sq ~�ή��q ~ q ~�9t 1142t 75pw        sq ~�ή�yq ~ q ~�9t 1142t 84pw@@�鹙�sq ~�ή�[q ~ q ~�9t 1143t 61pw        sq ~�ή�:q ~ q ~�9t 1143t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1144t 84pw@$      sq ~�ή��q ~ q ~�9t 1145t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1146t 75pw        sq ~�ή�}q ~ q ~�9t 1146t 84pw@5oz�G�sq ~�ή�_q ~ q ~�9t 1147t 61pw        sq ~�ή�>q ~ q ~�9t 1147t 84pw@$      sq ~�ή��q ~ q ~�9t 1148t 84pw@F�U�i�sq ~�ή�q ~ q ~�9t 1149t 75pw        sq ~�ή��q ~ q ~�9t 1149t 84pw@$      sq ~��Zw�0q ~ q ~�9t 115t 84pw@5oz�G�sq ~�ήVq ~ q ~�9t 1150t 84pw@@�鹙�sq ~�ήuq ~ q ~�9t 1151t 75pw        sq ~�ήq ~ q ~�9t 1151t 84pw@@�鹙�sq ~�ή
�q ~ q ~�9t 1152t 84pw@$      sq ~�ή�q ~ q ~�9t 1153t 61pw        sq ~�ή�q ~ q ~�9t 1153t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1154t 75pw        sq ~�ήZq ~ q ~�9t 1154t 84pw@@�鹙�sq ~�ήq ~ q ~�9t 1155t 84pw@@�鹙�sq ~�ή:q ~ q ~�9t 1156t 75pw        sq ~�ή�q ~ q ~�9t 1156t 84pw@@�鹙�sq ~�ή�q ~ q ~�9t 1157t 61pw        sq ~�ή�q ~ q ~�9t 1157t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1158t 75pw        sq ~�ή!^q ~ q ~�9t 1158t 84pw@@�鹙�sq ~�ή!}q ~ q ~�9t 1159t 75pw        sq ~�ή%q ~ q ~�9t 1159t 84pw@@�鹙�sq ~��Zw��q ~ q ~�9t 116t 84pw@5oz�G�sq ~�ήtq ~ q ~�9t 1160t 75pw        sq ~�ήw�q ~ q ~�9t 1160t 84pw@"D�^���sq ~�ήw�q ~ q ~�9t 1161t 75pw        sq ~�ή{vq ~ q ~�9t 1161t 84pw@F�U�i�sq ~�ή{�q ~ q ~�9t 1162t 75pw        sq ~�ή7q ~ q ~�9t 1162t 84pw@@�鹙�sq ~�ή{q ~ q ~�9t 1163t 61pw        sq ~�ή��q ~ q ~�9t 1163t 84pw@$      sq ~�ή~�q ~ q ~�9t 1164t 61pw        sq ~�ή��q ~ q ~�9t 1164t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1165t 61pw        sq ~�ή�zq ~ q ~�9t 1165t 84pw@5oz�G�sq ~�ή�\q ~ q ~�9t 1166t 61pw        sq ~�ή�;q ~ q ~�9t 1166t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1167t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1168t 61pw        sq ~�ή��q ~ q ~�9t 1168t 84pw@@�鹙�sq ~�ή�~q ~ q ~�9t 1169t 84pw@@�鹙�sq ~��Zwղq ~ q ~�9t 117t 84pw@$      sq ~�ή�5q ~ q ~�9t 1170t 61pw        sq ~�ή�q ~ q ~�9t 1170t 84pw@5oz�G�sq ~�ή�3q ~ q ~�9t 1171t 75pw        sq ~�ή��q ~ q ~�9t 1171t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1172t 75pw        sq ~�ή�q ~ q ~�9t 1172t 84pw@$      sq ~�ή�q ~ q ~�9t 1173t 75pw        sq ~�ή�Wq ~ q ~�9t 1173t 84pw@5oz�G�sq ~�ή�vq ~ q ~�9t 1174t 75pw        sq ~�ή�q ~ q ~�9t 1174t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1175t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1176t 61pw        sq ~�ή�q ~ q ~�9t 1176t 84pw@@�鹙�sq ~�ή�q ~ q ~�9t 1177t 75pw        sq ~�ή[q ~ q ~�9t 1177t 84pw@@�鹙�sq ~�ή=q ~ q ~�9t 1178t 61pw        sq ~�ή
q ~ q ~�9t 1178t 84pw@@�鹙�sq ~�ή
;q ~ q ~�9t 1179t 75pw        sq ~�ή�q ~ q ~�9t 1179t 84pw@5oz�G�sq ~��Zwєq ~ q ~�9t 118t 61pw        sq ~��Zw�sq ~ q ~�9t 118t 84pw@5oz�G�sq ~�ή\�q ~ q ~�9t 1180t 75pw        sq ~�ή`sq ~ q ~�9t 1180t 84pw@F�U�i�sq ~�ή\Uq ~ q ~�9t 1181t 61pw        sq ~�ήd4q ~ q ~�9t 1181t 84pw@@�鹙�sq ~�ή`q ~ q ~�9t 1182t 61pw        sq ~�ήg�q ~ q ~�9t 1182t 84pw@5oz�G�sq ~�ήhq ~ q ~�9t 1183t 75pw        sq ~�ήk�q ~ q ~�9t 1183t 84pw@5oz�G�sq ~�ήk�q ~ q ~�9t 1184t 75pw        sq ~�ήowq ~ q ~�9t 1184t 84pw@$      sq ~�ήkYq ~ q ~�9t 1185t 61pw        sq ~�ήs8q ~ q ~�9t 1185t 84pw@@�鹙�sq ~�ήv�q ~ q ~�9t 1186t 84pw@@�鹙�sq ~�ήz�q ~ q ~�9t 1187t 84pw@5oz�G�sq ~�ήv�q ~ q ~�9t 1188t 61pw        sq ~�ή~{q ~ q ~�9t 1188t 84pw@@�鹙�sq ~�ήz]q ~ q ~�9t 1189t 61pw        sq ~�ή�<q ~ q ~�9t 1189t 84pw@5oz�G�sq ~��Zwْq ~ q ~�9t 119t 75pw        sq ~��Zw�4q ~ q ~�9t 119t 84pw@$      sq ~�ή��q ~ q ~�9t 1190t 84pw@F�U�i�sq ~�ή��q ~ q ~�9t 1191t 75pw        sq ~�ήؓq ~ q ~�9t 1191t 84pw@5oz�G�sq ~�ή�uq ~ q ~�9t 1192t 61pw        sq ~�ή�Tq ~ q ~�9t 1192t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1193t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1194t 84pw@$      sq ~�ή��q ~ q ~�9t 1195t 75pw        sq ~�ή�q ~ q ~�9t 1195t 84pw@5oz�G�sq ~�ή�q ~ q ~�9t 1196t 75pw        sq ~�ή�Xq ~ q ~�9t 1196t 84pw@'�p��j�sq ~�ή�q ~ q ~�9t 1197t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1198t 61pw        sq ~�ή��q ~ q ~�9t 1198t 84pw@$      sq ~�ή�q ~ q ~�9t 1199t 61pw        sq ~�ή��q ~ q ~�9t 1199t 84pw@$      sq ~��W�(�q ~ q ~�9t 12t 13pw        sq ~��W�qq ~ q ~�9t 12t 4pw@$      sq ~��W�8�q ~ q ~�9t 12t 59pw@$      sq ~��Zx,(q ~ q ~�9t 120t 75pw        sq ~��Zx/�q ~ q ~�9t 120t 84pw@5oz�G�sq ~�ή"�Zq ~ q ~�9t 1200t 75pw        sq ~�ή"��q ~ q ~�9t 1200t 84pw@5oz�G�sq ~�ή"ؽq ~ q ~�9t 1201t 84pw@5oz�G�sq ~�ή"ԟq ~ q ~�9t 1202t 61pw        sq ~�ή"�~q ~ q ~�9t 1202t 84pw@@�鹙�sq ~�ή"�`q ~ q ~�9t 1203t 61pw        sq ~�ή"�?q ~ q ~�9t 1203t 84pw@$      sq ~�ή"�^q ~ q ~�9t 1204t 75pw        sq ~�ή"� q ~ q ~�9t 1204t 84pw@5oz�G�sq ~�ή"��q ~ q ~�9t 1205t 61pw        sq ~�ή"��q ~ q ~�9t 1205t 84pw@@�鹙�sq ~�ή"�q ~ q ~�9t 1206t 84pw@5oz�G�sq ~�ή"�Cq ~ q ~�9t 1207t 84pw@@�鹙�sq ~�ή"�bq ~ q ~�9t 1208t 75pw        sq ~�ή"�q ~ q ~�9t 1208t 84pw@5oz�G�sq ~�ή"�#q ~ q ~�9t 1209t 75pw        sq ~�ή"��q ~ q ~�9t 1209t 84pw@@�鹙�sq ~��Zx+�q ~ q ~�9t 121t 61pw        sq ~��Zx3�q ~ q ~�9t 121t 84pw@5oz�G�sq ~�ή#E�q ~ q ~�9t 1210t 75pw        sq ~�ή#I[q ~ q ~�9t 1210t 84pw@5oz�G�sq ~�ή#E=q ~ q ~�9t 1211t 61pw        sq ~�ή#Mq ~ q ~�9t 1211t 84pw@5oz�G�sq ~�ή#H�q ~ q ~�9t 1212t 61pw        sq ~�ή#P�q ~ q ~�9t 1212t 84pw@$      sq ~�ή#L�q ~ q ~�9t 1213t 61pw        sq ~�ή#T�q ~ q ~�9t 1213t 84pw@@�鹙�sq ~�ή#P�q ~ q ~�9t 1214t 61pw        sq ~�ή#X_q ~ q ~�9t 1214t 84pw@5oz�G�sq ~�ή#TAq ~ q ~�9t 1215t 61pw        sq ~�ή#\ q ~ q ~�9t 1215t 84pw@@�鹙�sq ~�ή#Xq ~ q ~�9t 1216t 61pw        sq ~�ή#_�q ~ q ~�9t 1216t 84pw@$      sq ~�ή#` q ~ q ~�9t 1217t 75pw        sq ~�ή#c�q ~ q ~�9t 1217t 84pw@@�鹙�sq ~�ή#c�q ~ q ~�9t 1218t 75pw        sq ~�ή#gcq ~ q ~�9t 1218t 84pw@$      sq ~�ή#cEq ~ q ~�9t 1219t 61pw        sq ~�ή#k$q ~ q ~�9t 1219t 84pw@F�U�i�sq ~��Zx/mq ~ q ~�9t 122t 61pw        sq ~��Zx7Lq ~ q ~�9t 122t 84pw@5oz�G�sq ~�ή#�q ~ q ~�9t 1220t 75pw        sq ~�ή#��q ~ q ~�9t 1220t 84pw@$      sq ~�ή#�{q ~ q ~�9t 1221t 84pw@5oz�G�sq ~�ή#�<q ~ q ~�9t 1222t 84pw@@�鹙�sq ~�ή#�[q ~ q ~�9t 1223t 75pw        sq ~�ή#��q ~ q ~�9t 1223t 84pw@5oz�G�sq ~�ή#̾q ~ q ~�9t 1224t 84pw@5oz�G�sq ~�ή#Ƞq ~ q ~�9t 1225t 61pw        sq ~�ή#�q ~ q ~�9t 1225t 84pw@@�鹙�sq ~�ή#Оq ~ q ~�9t 1226t 75pw        sq ~�ή#�@q ~ q ~�9t 1226t 84pw@F�U�i�sq ~�ή#�q ~ q ~�9t 1227t 84pw@5oz�G�sq ~�ή#� q ~ q ~�9t 1228t 75pw        sq ~�ή#��q ~ q ~�9t 1228t 84pw@$      sq ~�ή#��q ~ q ~�9t 1229t 75pw        sq ~�ή#߃q ~ q ~�9t 1229t 84pw@5oz�G�sq ~��Zx;q ~ q ~�9t 123t 84pw@@�鹙�sq ~�ή$.wq ~ q ~�9t 1230t 75pw        sq ~�ή$2q ~ q ~�9t 1230t 84pw@@�鹙�sq ~�ή$-�q ~ q ~�9t 1231t 61pw        sq ~�ή$5�q ~ q ~�9t 1231t 84pw@@�鹙�sq ~�ή$5�q ~ q ~�9t 1232t 75pw        sq ~�ή$9�q ~ q ~�9t 1232t 84pw@5oz�G�sq ~�ή$=\q ~ q ~�9t 1233t 84pw@5oz�G�sq ~�ή$Aq ~ q ~�9t 1234t 84pw@$      sq ~�ή$<�q ~ q ~�9t 1235t 61pw        sq ~�ή$D�q ~ q ~�9t 1235t 84pw@5oz�G�sq ~�ή$@�q ~ q ~�9t 1236t 61pw        sq ~�ή$H�q ~ q ~�9t 1236t 84pw@@�鹙�sq ~�ή$L`q ~ q ~�9t 1237t 84pw@5oz�G�sq ~�ή$Lq ~ q ~�9t 1238t 75pw        sq ~�ή$P!q ~ q ~�9t 1238t 84pw@M]��%��sq ~�ή$Lq ~ q ~�9t 1239t 61pw        sq ~�ή$S�q ~ q ~�9t 1239t 84pw@5oz�G�sq ~��Zx>�q ~ q ~�9t 124t 84pw@@�鹙�sq ~�ή$�xq ~ q ~�9t 1240t 84pw@$      sq ~�ή$�9q ~ q ~�9t 1241t 84pw@#�׭�Bsq ~�ή$��q ~ q ~�9t 1242t 84pw@$      sq ~�ή$��q ~ q ~�9t 1243t 84pw@5oz�G�sq ~�ή$�|q ~ q ~�9t 1244t 84pw@5oz�G�sq ~�ή$��q ~ q ~�9t 1245t 75pw        sq ~�ή$�=q ~ q ~�9t 1245t 84pw@5oz�G�sq ~�ή$�\q ~ q ~�9t 1246t 75pw        sq ~�ή$��q ~ q ~�9t 1246t 84pw@5oz�G�sq ~�ή$�q ~ q ~�9t 1247t 75pw        sq ~�ή$��q ~ q ~�9t 1247t 84pw@5oz�G�sq ~�ή$Āq ~ q ~�9t 1248t 84pw@$      sq ~�ή$�Aq ~ q ~�9t 1249t 84pw@5oz�G�sq ~��Zx:�q ~ q ~�9t 125t 61pw        sq ~��ZxB�q ~ q ~�9t 125t 84pw@$      sq ~�ή%5q ~ q ~�9t 1250t 75pw        sq ~�ή%�q ~ q ~�9t 1250t 84pw@5oz�G�sq ~�ή%�q ~ q ~�9t 1251t 75pw        sq ~�ή%�q ~ q ~�9t 1251t 84pw@5oz�G�sq ~�ή%�q ~ q ~�9t 1252t 75pw        sq ~�ή%"Yq ~ q ~�9t 1252t 84pw@5oz�G�sq ~�ή%"xq ~ q ~�9t 1253t 75pw        sq ~�ή%&q ~ q ~�9t 1253t 84pw@@�鹙�sq ~�ή%!�q ~ q ~�9t 1254t 61pw        sq ~�ή%)�q ~ q ~�9t 1254t 84pw@@�鹙�sq ~�ή%-�q ~ q ~�9t 1255t 84pw@@�鹙�sq ~�ή%-�q ~ q ~�9t 1256t 75pw        sq ~�ή%1]q ~ q ~�9t 1256t 84pw@$      sq ~�ή%-?q ~ q ~�9t 1257t 61pw        sq ~�ή%5q ~ q ~�9t 1257t 84pw@5	H�>sq ~�ή%1 q ~ q ~�9t 1258t 61pw        sq ~�ή%8�q ~ q ~�9t 1258t 84pw@#�����Jsq ~�ή%4�q ~ q ~�9t 1259t 61pw        sq ~�ή%<�q ~ q ~�9t 1259t 84pw@$      sq ~��ZxB�q ~ q ~�9t 126t 75pw        sq ~��ZxFPq ~ q ~�9t 126t 84pw@@�鹙�sq ~�ή%��q ~ q ~�9t 1260t 75pw        sq ~�ή%�6q ~ q ~�9t 1260t 84pw@@�鹙�sq ~�ή%��q ~ q ~�9t 1261t 84pw@$      sq ~�ή%��q ~ q ~�9t 1262t 84pw@5oz�G�sq ~�ή%��q ~ q ~�9t 1263t 75pw        sq ~�ή%�yq ~ q ~�9t 1263t 84pw@@�鹙�sq ~�ή%��q ~ q ~�9t 1264t 75pw        sq ~�ή%�:q ~ q ~�9t 1264t 84pw@$      sq ~�ή%�Yq ~ q ~�9t 1265t 75pw        sq ~�ή%��q ~ q ~�9t 1265t 84pw@5oz�G�sq ~�ή%�q ~ q ~�9t 1266t 75pw        sq ~�ή%��q ~ q ~�9t 1266t 84pw@$      sq ~�ή%��q ~ q ~�9t 1267t 61pw        sq ~�ή%�}q ~ q ~�9t 1267t 84pw@$      sq ~�ή%�_q ~ q ~�9t 1268t 61pw        sq ~�ή%�>q ~ q ~�9t 1268t 84pw@5oz�G�sq ~�ή%��q ~ q ~�9t 1269t 84pw@5oz�G�sq ~��ZxB2q ~ q ~�9t 127t 61pw        sq ~��ZxJq ~ q ~�9t 127t 84pw@$      sq ~�ή%��q ~ q ~�9t 1270t 75pw        sq ~�ή&�q ~ q ~�9t 1270t 84pw@@�鹙�sq ~�ή&Vq ~ q ~�9t 1271t 84pw@5oz�G�sq ~�ή&uq ~ q ~�9t 1272t 75pw        sq ~�ή&q ~ q ~�9t 1272t 84pw@$      sq ~�ή&�q ~ q ~�9t 1273t 61pw        sq ~�ή&�q ~ q ~�9t 1273t 84pw@5oz�G�sq ~�ή&�q ~ q ~�9t 1274t 84pw@F�U�i�sq ~�ή&Zq ~ q ~�9t 1275t 84pw@@�鹙�sq ~�ή&yq ~ q ~�9t 1276t 75pw        sq ~�ή&q ~ q ~�9t 1276t 84pw@@�鹙�sq ~�ή&�q ~ q ~�9t 1277t 61pw        sq ~�ή&�q ~ q ~�9t 1277t 84pw@$      sq ~�ή&!�q ~ q ~�9t 1278t 84pw@+�,W8�*sq ~�ή&!�q ~ q ~�9t 1279t 75pw        sq ~�ή&%^q ~ q ~�9t 1279t 84pw@5oz�G�sq ~��ZxM�q ~ q ~�9t 128t 84pw@@�鹙�sq ~�ή&pq ~ q ~�9t 1280t 61pw        sq ~�ή&w�q ~ q ~�9t 1280t 84pw@@�鹙�sq ~�ή&{�q ~ q ~�9t 1281t 84pw@@�鹙�sq ~�ή&w�q ~ q ~�9t 1282t 61pw        sq ~�ή&vq ~ q ~�9t 1282t 84pw@$      sq ~�ή&�q ~ q ~�9t 1283t 75pw        sq ~�ή&�7q ~ q ~�9t 1283t 84pw@$      sq ~�ή&q ~ q ~�9t 1284t 61pw        sq ~�ή&��q ~ q ~�9t 1284t 84pw@@�鹙�sq ~�ή&�q ~ q ~�9t 1285t 75pw        sq ~�ή&��q ~ q ~�9t 1285t 84pw@5oz�G�sq ~�ή&��q ~ q ~�9t 1286t 75pw        sq ~�ή&�zq ~ q ~�9t 1286t 84pw@@�鹙�sq ~�ή&��q ~ q ~�9t 1287t 75pw        sq ~�ή&�;q ~ q ~�9t 1287t 84pw@5oz�G�sq ~�ή&��q ~ q ~�9t 1288t 84pw@5oz�G�sq ~�ή&��q ~ q ~�9t 1289t 61pw        sq ~�ή&��q ~ q ~�9t 1289t 84pw@5oz�G�sq ~��ZxI�q ~ q ~�9t 129t 61pw        sq ~��ZxQ�q ~ q ~�9t 129t 84pw@5oz�G�sq ~�ή&�tq ~ q ~�9t 1290t 61pw        sq ~�ή&�Sq ~ q ~�9t 1290t 84pw@5oz�G�sq ~�ή&�rq ~ q ~�9t 1291t 75pw        sq ~�ή&�q ~ q ~�9t 1291t 84pw@@�鹙�sq ~�ή&��q ~ q ~�9t 1292t 61pw        sq ~�ή&��q ~ q ~�9t 1292t 84pw@$      sq ~�ή&��q ~ q ~�9t 1293t 84pw@@�鹙�sq ~�ή&�Wq ~ q ~�9t 1294t 84pw@$      sq ~�ή&�vq ~ q ~�9t 1295t 75pw        sq ~�ή&�q ~ q ~�9t 1295t 84pw@5oz�G�sq ~�ή'�q ~ q ~�9t 1296t 84pw@5oz�G�sq ~�ή&��q ~ q ~�9t 1297t 61pw        sq ~�ή'�q ~ q ~�9t 1297t 84pw@5oz�G�sq ~�ή'|q ~ q ~�9t 1298t 61pw        sq ~�ή'
[q ~ q ~�9t 1298t 84pw@5oz�G�sq ~�ή'
zq ~ q ~�9t 1299t 75pw        sq ~�ή'q ~ q ~�9t 1299t 84pw@5oz�G�sq ~��W�,�q ~ q ~�9t 13t 14pw        sq ~��W�,�q ~ q ~�9t 13t 15pw���܅ib?sq ~��W�7�q ~ q ~�9t 13t 43pw@$      sq ~��Zx��q ~ q ~�9t 130t 75pw        sq ~��Zx�)q ~ q ~�9t 130t 84pw@@�鹙�sq ~�ή0��q ~ q ~�9t 1300t 75pw        sq ~�ή0�}q ~ q ~�9t 1300t 84pw@$      sq ~�ή0�>q ~ q ~�9t 1301t 84pw@@�鹙�sq ~�ή0�]q ~ q ~�9t 1302t 75pw        sq ~�ή0��q ~ q ~�9t 1302t 84pw@@�鹙�sq ~�ή0�q ~ q ~�9t 1303t 75pw        sq ~�ή0��q ~ q ~�9t 1303t 84pw@$      sq ~�ή0��q ~ q ~�9t 1304t 84pw@5oz�G�sq ~�ή0�Bq ~ q ~�9t 1305t 84pw@5oz�G�sq ~�ή1q ~ q ~�9t 1306t 84pw@5oz�G�sq ~�ή1�q ~ q ~�9t 1307t 84pw@M]��%��sq ~�ή1�q ~ q ~�9t 1308t 61pw        sq ~�ή1
�q ~ q ~�9t 1308t 84pw@@�鹙�sq ~�ή1
�q ~ q ~�9t 1309t 75pw        sq ~�ή1Fq ~ q ~�9t 1309t 84pw@5oz�G�sq ~��Zx�Hq ~ q ~�9t 131t 75pw        sq ~��Zx��q ~ q ~�9t 131t 84pw@$      sq ~�ή1`�q ~ q ~�9t 1310t 84pw@@�鹙�sq ~�ή1\�q ~ q ~�9t 1311t 61pw        sq ~�ή1d�q ~ q ~�9t 1311t 84pw@$      sq ~�ή1h^q ~ q ~�9t 1312t 84pw@5oz�G�sq ~�ή1d@q ~ q ~�9t 1313t 61pw        sq ~�ή1lq ~ q ~�9t 1313t 84pw@5oz�G�sq ~�ή1o�q ~ q ~�9t 1314t 84pw@5oz�G�sq ~�ή1k�q ~ q ~�9t 1315t 61pw        sq ~�ή1s�q ~ q ~�9t 1315t 84pw@$      sq ~�ή1wbq ~ q ~�9t 1316t 84pw@@�鹙�sq ~�ή1w�q ~ q ~�9t 1317t 75pw        sq ~�ή1{#q ~ q ~�9t 1317t 84pw@M]��%��sq ~�ή1wq ~ q ~�9t 1318t 61pw        sq ~�ή1~�q ~ q ~�9t 1318t 84pw@$      sq ~�ή1z�q ~ q ~�9t 1319t 61pw        sq ~�ή1��q ~ q ~�9t 1319t 84pw@F�U�i�sq ~��Zx��q ~ q ~�9t 132t 61pw        sq ~��Zx��q ~ q ~�9t 132t 84pw@5oz�G�sq ~�ή1�\q ~ q ~�9t 1320t 61pw        sq ~�ή1�;q ~ q ~�9t 1320t 84pw@5oz�G�sq ~�ή1��q ~ q ~�9t 1321t 84pw@@�鹙�sq ~�ή1��q ~ q ~�9t 1322t 61pw        sq ~�ή1ܽq ~ q ~�9t 1322t 84pw@$      sq ~�ή1��q ~ q ~�9t 1323t 75pw        sq ~�ή1�~q ~ q ~�9t 1323t 84pw@F�U�i�sq ~�ή1��q ~ q ~�9t 1324t 75pw        sq ~�ή1�?q ~ q ~�9t 1324t 84pw@5oz�G�sq ~�ή1� q ~ q ~�9t 1325t 84pw@@�鹙�sq ~�ή1��q ~ q ~�9t 1326t 61pw        sq ~�ή1��q ~ q ~�9t 1326t 84pw@5oz�G�sq ~�ή1�q ~ q ~�9t 1327t 84pw@$      sq ~�ή1�dq ~ q ~�9t 1328t 61pw        sq ~�ή1�Cq ~ q ~�9t 1328t 84pw@$      sq ~�ή1�%q ~ q ~�9t 1329t 61pw        sq ~�ή1�q ~ q ~�9t 1329t 84pw@$      sq ~��Zx��q ~ q ~�9t 133t 75pw        sq ~��Zx�lq ~ q ~�9t 133t 84pw@@�鹙�sq ~�ή2A�q ~ q ~�9t 1330t 61pw        sq ~�ή2I�q ~ q ~�9t 1330t 84pw@5oz�G�sq ~�ή2M[q ~ q ~�9t 1331t 84pw@@�鹙�sq ~�ή2Mzq ~ q ~�9t 1332t 75pw        sq ~�ή2Qq ~ q ~�9t 1332t 84pw@5oz�G�sq ~�ή2T�q ~ q ~�9t 1333t 84pw@@�鹙�sq ~�ή2T�q ~ q ~�9t 1334t 75pw        sq ~�ή2X�q ~ q ~�9t 1334t 84pw@7�ÓHrsq ~�ή2X�q ~ q ~�9t 1335t 75pw        sq ~�ή2\_q ~ q ~�9t 1335t 84pw@5oz�G�sq ~�ή2` q ~ q ~�9t 1336t 84pw@$      sq ~�ή2c�q ~ q ~�9t 1337t 84pw@@�鹙�sq ~�ή2d q ~ q ~�9t 1338t 75pw        sq ~�ή2g�q ~ q ~�9t 1338t 84pw@5oz�G�sq ~�ή2c�q ~ q ~�9t 1339t 61pw        sq ~�ή2kcq ~ q ~�9t 1339t 84pw@5oz�G�sq ~��Zx��q ~ q ~�9t 134t 75pw        sq ~��Zx�-q ~ q ~�9t 134t 84pw@$      sq ~�ή2�Wq ~ q ~�9t 1340t 75pw        sq ~�ή2��q ~ q ~�9t 1340t 84pw@@�鹙�sq ~�ή2��q ~ q ~�9t 1341t 84pw@%����i%sq ~�ή2��q ~ q ~�9t 1342t 61pw        sq ~�ή2�{q ~ q ~�9t 1342t 84pw@$      sq ~�ή2�<q ~ q ~�9t 1343t 84pw@$      sq ~�ή2�[q ~ q ~�9t 1344t 75pw        sq ~�ή2��q ~ q ~�9t 1344t 84pw@@�鹙�sq ~�ή2оq ~ q ~�9t 1345t 84pw@5oz�G�sq ~�ή2̠q ~ q ~�9t 1346t 61pw        sq ~�ή2�q ~ q ~�9t 1346t 84pw@$      sq ~�ή2�aq ~ q ~�9t 1347t 61pw        sq ~�ή2�@q ~ q ~�9t 1347t 84pw@5oz�G�sq ~�ή2�"q ~ q ~�9t 1348t 61pw        sq ~�ή2�q ~ q ~�9t 1348t 84pw@$      sq ~�ή2� q ~ q ~�9t 1349t 75pw        sq ~�ή2��q ~ q ~�9t 1349t 84pw@@�鹙�sq ~��Zx�q ~ q ~�9t 135t 61pw        sq ~��Zx��q ~ q ~�9t 135t 84pw@$      sq ~�ή3*yq ~ q ~�9t 1350t 61pw        sq ~�ή32Xq ~ q ~�9t 1350t 84pw@$      sq ~�ή3.:q ~ q ~�9t 1351t 61pw        sq ~�ή36q ~ q ~�9t 1351t 84pw@$      sq ~�ή31�q ~ q ~�9t 1352t 61pw        sq ~�ή39�q ~ q ~�9t 1352t 84pw@$      sq ~�ή39�q ~ q ~�9t 1353t 75pw        sq ~�ή3=�q ~ q ~�9t 1353t 84pw@$      sq ~�ή3A\q ~ q ~�9t 1354t 84pw@$      sq ~�ή3Eq ~ q ~�9t 1355t 84pw@5oz�G�sq ~�ή3@�q ~ q ~�9t 1356t 61pw        sq ~�ή3H�q ~ q ~�9t 1356t 84pw@5oz�G�sq ~�ή3H�q ~ q ~�9t 1357t 75pw        sq ~�ή3L�q ~ q ~�9t 1357t 84pw@@�鹙�sq ~�ή3L�q ~ q ~�9t 1358t 75pw        sq ~�ή3P`q ~ q ~�9t 1358t 84pw@5oz�G�sq ~�ή3T!q ~ q ~�9t 1359t 84pw@$      sq ~��Zx�q ~ q ~�9t 136t 75pw        sq ~��Zx��q ~ q ~�9t 136t 84pw@@�鹙�sq ~�ή3�q ~ q ~�9t 1360t 75pw        sq ~�ή3��q ~ q ~�9t 1360t 84pw@5oz�G�sq ~�ή3��q ~ q ~�9t 1361t 75pw        sq ~�ή3�xq ~ q ~�9t 1361t 84pw@5oz�G�sq ~�ή3�Zq ~ q ~�9t 1362t 61pw        sq ~�ή3�9q ~ q ~�9t 1362t 84pw@$      sq ~�ή3�Xq ~ q ~�9t 1363t 75pw        sq ~�ή3��q ~ q ~�9t 1363t 84pw@5oz�G�sq ~�ή3��q ~ q ~�9t 1364t 61pw        sq ~�ή3��q ~ q ~�9t 1364t 84pw@$      sq ~�ή3�|q ~ q ~�9t 1365t 84pw@5oz�G�sq ~�ή3�^q ~ q ~�9t 1366t 61pw        sq ~�ή3�=q ~ q ~�9t 1366t 84pw@%���L_sq ~�ή3�\q ~ q ~�9t 1367t 75pw        sq ~�ή3��q ~ q ~�9t 1367t 84pw@@�鹙�sq ~�ή3�q ~ q ~�9t 1368t 75pw        sq ~�ή3Ŀq ~ q ~�9t 1368t 84pw@5oz�G�sq ~�ή3��q ~ q ~�9t 1369t 61pw        sq ~�ή3Ȁq ~ q ~�9t 1369t 84pw@$      sq ~��Zx�pq ~ q ~�9t 137t 84pw@5oz�G�sq ~�ή47q ~ q ~�9t 1370t 61pw        sq ~�ή4q ~ q ~�9t 1370t 84pw@$      sq ~�ή45q ~ q ~�9t 1371t 75pw        sq ~�ή4�q ~ q ~�9t 1371t 84pw@5oz�G�sq ~�ή4"�q ~ q ~�9t 1372t 84pw@$      sq ~�ή4"�q ~ q ~�9t 1373t 75pw        sq ~�ή4&Yq ~ q ~�9t 1373t 84pw@$      sq ~�ή4&xq ~ q ~�9t 1374t 75pw        sq ~�ή4*q ~ q ~�9t 1374t 84pw@5oz�G�sq ~�ή4*9q ~ q ~�9t 1375t 75pw        sq ~�ή4-�q ~ q ~�9t 1375t 84pw@F�U�i�sq ~�ή41�q ~ q ~�9t 1376t 84pw@@�鹙�sq ~�ή4-~q ~ q ~�9t 1377t 61pw        sq ~�ή45]q ~ q ~�9t 1377t 84pw@5oz�G�sq ~�ή45|q ~ q ~�9t 1378t 75pw        sq ~�ή49q ~ q ~�9t 1378t 84pw@5oz�G�sq ~�ή4<�q ~ q ~�9t 1379t 84pw@$      sq ~��Zx�1q ~ q ~�9t 138t 84pw@5oz�G�sq ~�ή4�uq ~ q ~�9t 1380t 84pw@$      sq ~�ή4��q ~ q ~�9t 1381t 75pw        sq ~�ή4�6q ~ q ~�9t 1381t 84pw@$      sq ~�ή4�q ~ q ~�9t 1382t 61pw        sq ~�ή4��q ~ q ~�9t 1382t 84pw@@�鹙�sq ~�ή4�q ~ q ~�9t 1383t 75pw        sq ~�ή4��q ~ q ~�9t 1383t 84pw@5oz�G�sq ~�ή4��q ~ q ~�9t 1384t 61pw        sq ~�ή4�yq ~ q ~�9t 1384t 84pw@F�U�i�sq ~�ή4��q ~ q ~�9t 1385t 75pw        sq ~�ή4�:q ~ q ~�9t 1385t 84pw@$      sq ~�ή4�q ~ q ~�9t 1386t 61pw        sq ~�ή4��q ~ q ~�9t 1386t 84pw@@�鹙�sq ~�ή4��q ~ q ~�9t 1387t 84pw@@�鹙�sq ~�ή4��q ~ q ~�9t 1388t 75pw        sq ~�ή4�}q ~ q ~�9t 1388t 84pw@5oz�G�sq ~�ή4�_q ~ q ~�9t 1389t 61pw        sq ~�ή4�>q ~ q ~�9t 1389t 84pw@@�鹙�sq ~��Zx��q ~ q ~�9t 139t 84pw@@�鹙�sq ~�ή4��q ~ q ~�9t 1390t 61pw        sq ~�ή5�q ~ q ~�9t 1390t 84pw@@�鹙�sq ~�ή5�q ~ q ~�9t 1391t 84pw@F�U�i�sq ~�ή5�q ~ q ~�9t 1392t 75pw        sq ~�ή5Vq ~ q ~�9t 1392t 84pw@$      sq ~�ή58q ~ q ~�9t 1393t 61pw        sq ~�ή5q ~ q ~�9t 1393t 84pw@F�U�i�sq ~�ή5�q ~ q ~�9t 1394t 84pw@@�鹙�sq ~�ή5�q ~ q ~�9t 1395t 61pw        sq ~�ή5�q ~ q ~�9t 1395t 84pw@$      sq ~�ή5�q ~ q ~�9t 1396t 75pw        sq ~�ή5Zq ~ q ~�9t 1396t 84pw@$      sq ~�ή5<q ~ q ~�9t 1397t 61pw        sq ~�ή5q ~ q ~�9t 1397t 84pw@$      sq ~�ή5:q ~ q ~�9t 1398t 75pw        sq ~�ή5!�q ~ q ~�9t 1398t 84pw@5oz�G�sq ~�ή5%�q ~ q ~�9t 1399t 84pw@%�����sq ~��W�0�q ~ q ~�9t 14t 16pw        sq ~��W�>�q ~ q ~�9t 14t 50pw        sq ~��W�x�q ~ q ~�9t 14t 6pw@$      sq ~��Zy�q ~ q ~�9t 140t 61pw        sq ~��Zy�q ~ q ~�9t 140t 84pw@@�鹙�sq ~�ή? \q ~ q ~�9t 1400t 75pw        sq ~�ή?�q ~ q ~�9t 1400t 84pw@5oz�G�sq ~�ή>��q ~ q ~�9t 1401t 61pw        sq ~�ή?�q ~ q ~�9t 1401t 84pw@$      sq ~�ή?�q ~ q ~�9t 1402t 84pw@$      sq ~�ή?�q ~ q ~�9t 1403t 75pw        sq ~�ή?Aq ~ q ~�9t 1403t 84pw@5oz�G�sq ~�ή?`q ~ q ~�9t 1404t 75pw        sq ~�ή?q ~ q ~�9t 1404t 84pw@$      sq ~�ή?!q ~ q ~�9t 1405t 75pw        sq ~�ή?�q ~ q ~�9t 1405t 84pw@@�鹙�sq ~�ή?�q ~ q ~�9t 1406t 75pw        sq ~�ή?�q ~ q ~�9t 1406t 84pw@@�鹙�sq ~�ή?fq ~ q ~�9t 1407t 61pw        sq ~�ή?Eq ~ q ~�9t 1407t 84pw@@�鹙�sq ~�ή?'q ~ q ~�9t 1408t 61pw        sq ~�ή?"q ~ q ~�9t 1408t 84pw@$      sq ~�ή?�q ~ q ~�9t 1409t 61pw        sq ~�ή?%�q ~ q ~�9t 1409t 84pw@$      sq ~��Zyjq ~ q ~�9t 141t 61pw        sq ~��ZyIq ~ q ~�9t 141t 84pw@5oz�G�sq ~�ή?x]q ~ q ~�9t 1410t 84pw@5oz�G�sq ~�ή?|q ~ q ~�9t 1411t 84pw@6eeÐGpsq ~�ή?�q ~ q ~�9t 1412t 84pw@$      sq ~�ή?��q ~ q ~�9t 1413t 84pw@@�鹙�sq ~�ή?�aq ~ q ~�9t 1414t 84pw@@�鹙�sq ~�ή?�Cq ~ q ~�9t 1415t 61pw        sq ~�ή?�"q ~ q ~�9t 1415t 84pw@F�U�i�sq ~�ή?�q ~ q ~�9t 1416t 61pw        sq ~�ή?��q ~ q ~�9t 1416t 84pw@@�鹙�sq ~�ή?�q ~ q ~�9t 1417t 75pw        sq ~�ή?��q ~ q ~�9t 1417t 84pw@5oz�G�sq ~�ή?��q ~ q ~�9t 1418t 61pw        sq ~�ή?�eq ~ q ~�9t 1418t 84pw@@�鹙�sq ~�ή?��q ~ q ~�9t 1419t 75pw        sq ~�ή?�&q ~ q ~�9t 1419t 84pw@@�鹙�sq ~��Zy 
q ~ q ~�9t 142t 84pw@$      sq ~�ή?��q ~ q ~�9t 1420t 61pw        sq ~�ή?�q ~ q ~�9t 1420t 84pw@5oz�G�sq ~�ή?�q ~ q ~�9t 1421t 61pw        sq ~�ή?�}q ~ q ~�9t 1421t 84pw@$      sq ~�ή?�_q ~ q ~�9t 1422t 61pw        sq ~�ή?�>q ~ q ~�9t 1422t 84pw@@�鹙�sq ~�ή?� q ~ q ~�9t 1423t 61pw        sq ~�ή?��q ~ q ~�9t 1423t 84pw@$      sq ~�ή?�q ~ q ~�9t 1424t 75pw        sq ~�ή?��q ~ q ~�9t 1424t 84pw@5oz�G�sq ~�ή?��q ~ q ~�9t 1425t 61pw        sq ~�ή?��q ~ q ~�9t 1425t 84pw@$      sq ~�ή?�cq ~ q ~�9t 1426t 61pw        sq ~�ή@Bq ~ q ~�9t 1426t 84pw@@�鹙�sq ~�ή?�$q ~ q ~�9t 1427t 61pw        sq ~�ή@q ~ q ~�9t 1427t 84pw@$      sq ~�ή@
�q ~ q ~�9t 1428t 84pw@5oz�G�sq ~�ή@�q ~ q ~�9t 1429t 84pw@$      sq ~��Zy )q ~ q ~�9t 143t 75pw        sq ~��Zy#�q ~ q ~�9t 143t 84pw@5oz�G�sq ~�ή@Y<q ~ q ~�9t 1430t 61pw        sq ~�ή@aq ~ q ~�9t 1430t 84pw@5oz�G�sq ~�ή@\�q ~ q ~�9t 1431t 61pw        sq ~�ή@d�q ~ q ~�9t 1431t 84pw@@�鹙�sq ~�ή@d�q ~ q ~�9t 1432t 75pw        sq ~�ή@h�q ~ q ~�9t 1432t 84pw@5oz�G�sq ~�ή@l^q ~ q ~�9t 1433t 84pw@5oz�G�sq ~�ή@l}q ~ q ~�9t 1434t 75pw        sq ~�ή@pq ~ q ~�9t 1434t 84pw@F�U�i�sq ~�ή@lq ~ q ~�9t 1435t 61pw        sq ~�ή@s�q ~ q ~�9t 1435t 84pw@@�鹙�sq ~�ή@o�q ~ q ~�9t 1436t 61pw        sq ~�ή@w�q ~ q ~�9t 1436t 84pw@$      sq ~�ή@s�q ~ q ~�9t 1437t 61pw        sq ~�ή@{bq ~ q ~�9t 1437t 84pw@@�鹙�sq ~�ή@{�q ~ q ~�9t 1438t 75pw        sq ~�ή@#q ~ q ~�9t 1438t 84pw@@�鹙�sq ~�ή@��q ~ q ~�9t 1439t 84pw@$      sq ~��Zy'�q ~ q ~�9t 144t 84pw@F�U�i�sq ~�ή@��q ~ q ~�9t 1440t 75pw        sq ~�ή@�zq ~ q ~�9t 1440t 84pw@5oz�G�sq ~�ή@ՙq ~ q ~�9t 1441t 75pw        sq ~�ή@�;q ~ q ~�9t 1441t 84pw@5oz�G�sq ~�ή@��q ~ q ~�9t 1442t 84pw@5oz�G�sq ~�ή@�q ~ q ~�9t 1443t 75pw        sq ~�ή@�q ~ q ~�9t 1443t 84pw@@�鹙�sq ~�ή@��q ~ q ~�9t 1444t 75pw        sq ~�ή@�~q ~ q ~�9t 1444t 84pw@5oz�G�sq ~�ή@�q ~ q ~�9t 1445t 75pw        sq ~�ή@�?q ~ q ~�9t 1445t 84pw@@�鹙�sq ~�ή@� q ~ q ~�9t 1446t 84pw@$>g�	��sq ~�ή@��q ~ q ~�9t 1447t 61pw        sq ~�ή@��q ~ q ~�9t 1447t 84pw@5oz�G�sq ~�ή@��q ~ q ~�9t 1448t 75pw        sq ~�ή@�q ~ q ~�9t 1448t 84pw@5oz�G�sq ~�ή@�q ~ q ~�9t 1449t 75pw        sq ~�ή@�Cq ~ q ~�9t 1449t 84pw@$      sq ~��Zy#nq ~ q ~�9t 145t 61pw        sq ~��Zy+Mq ~ q ~�9t 145t 84pw@5oz�G�sq ~�ήAF7q ~ q ~�9t 1450t 75pw        sq ~�ήAI�q ~ q ~�9t 1450t 84pw@@�鹙�sq ~�ήAI�q ~ q ~�9t 1451t 75pw        sq ~�ήAM�q ~ q ~�9t 1451t 84pw@5oz�G�sq ~�ήAI|q ~ q ~�9t 1452t 61pw        sq ~�ήAQ[q ~ q ~�9t 1452t 84pw@5oz�G�sq ~�ήAUq ~ q ~�9t 1453t 84pw@5oz�G�sq ~�ήAX�q ~ q ~�9t 1454t 84pw@$      sq ~�ήAT�q ~ q ~�9t 1455t 61pw        sq ~�ήA\�q ~ q ~�9t 1455t 84pw@5oz�G�sq ~�ήA`_q ~ q ~�9t 1456t 84pw@5oz�G�sq ~�ήA\Aq ~ q ~�9t 1457t 61pw        sq ~�ήAd q ~ q ~�9t 1457t 84pw@5oz�G�sq ~�ήAd?q ~ q ~�9t 1458t 75pw        sq ~�ήAg�q ~ q ~�9t 1458t 84pw@$      sq ~�ήAc�q ~ q ~�9t 1459t 61pw        sq ~�ήAk�q ~ q ~�9t 1459t 84pw@@�鹙�sq ~��Zy+lq ~ q ~�9t 146t 75pw        sq ~��Zy/q ~ q ~�9t 146t 84pw@@�鹙�sq ~�ήA�8q ~ q ~�9t 1460t 84pw@F�U�i�sq ~�ήA�Wq ~ q ~�9t 1461t 75pw        sq ~�ήA��q ~ q ~�9t 1461t 84pw@$      sq ~�ήAźq ~ q ~�9t 1462t 84pw@5oz�G�sq ~�ήA�{q ~ q ~�9t 1463t 84pw@5oz�G�sq ~�ήA�<q ~ q ~�9t 1464t 84pw@5oz�G�sq ~�ήA��q ~ q ~�9t 1465t 84pw@@�鹙�sq ~�ήAԾq ~ q ~�9t 1466t 84pw@$      sq ~�ήA��q ~ q ~�9t 1467t 75pw        sq ~�ήA�q ~ q ~�9t 1467t 84pw@&      sq ~�ήA�@q ~ q ~�9t 1468t 84pw@@�鹙�sq ~�ήA�"q ~ q ~�9t 1469t 61pw        sq ~�ήA�q ~ q ~�9t 1469t 84pw@5oz�G�sq ~��Zy2�q ~ q ~�9t 147t 84pw@$      sq ~�ήB*�q ~ q ~�9t 1470t 61pw        sq ~�ήB2�q ~ q ~�9t 1470t 84pw@@�鹙�sq ~�ήB6Xq ~ q ~�9t 1471t 84pw@@�鹙�sq ~�ήB2:q ~ q ~�9t 1472t 61pw        sq ~�ήB:q ~ q ~�9t 1472t 84pw@$      sq ~�ήB5�q ~ q ~�9t 1473t 61pw        sq ~�ήB=�q ~ q ~�9t 1473t 84pw@@�鹙�sq ~�ήB=�q ~ q ~�9t 1474t 75pw        sq ~�ήBA�q ~ q ~�9t 1474t 84pw@$      sq ~�ήBE\q ~ q ~�9t 1475t 84pw@@�鹙�sq ~�ήBE{q ~ q ~�9t 1476t 75pw        sq ~�ήBIq ~ q ~�9t 1476t 84pw@$      sq ~�ήBL�q ~ q ~�9t 1477t 84pw@5oz�G�sq ~�ήBL�q ~ q ~�9t 1478t 75pw        sq ~�ήBP�q ~ q ~�9t 1478t 84pw@F�U�i�sq ~�ήBP�q ~ q ~�9t 1479t 75pw        sq ~�ήBT`q ~ q ~�9t 1479t 84pw@@�鹙�sq ~��Zy6�q ~ q ~�9t 148t 84pw@$      sq ~�ήB�Tq ~ q ~�9t 1480t 75pw        sq ~�ήB��q ~ q ~�9t 1480t 84pw@@�鹙�sq ~�ήB��q ~ q ~�9t 1481t 84pw@5oz�G�sq ~�ήB��q ~ q ~�9t 1482t 61pw        sq ~�ήB�xq ~ q ~�9t 1482t 84pw@5oz�G�sq ~�ήB�9q ~ q ~�9t 1483t 84pw@$      sq ~�ήB�q ~ q ~�9t 1484t 61pw        sq ~�ήB��q ~ q ~�9t 1484t 84pw@5oz�G�sq ~�ήB�q ~ q ~�9t 1485t 75pw        sq ~�ήB��q ~ q ~�9t 1485t 84pw@@�鹙�sq ~�ήB��q ~ q ~�9t 1486t 61pw        sq ~�ήB�|q ~ q ~�9t 1486t 84pw@5oz�G�sq ~�ήB�=q ~ q ~�9t 1487t 84pw@5oz�G�sq ~�ήB��q ~ q ~�9t 1488t 84pw@5oz�G�sq ~�ήBȿq ~ q ~�9t 1489t 84pw@5oz�G�sq ~��Zy:Qq ~ q ~�9t 149t 84pw@'��D�;^sq ~�ήC�q ~ q ~�9t 1490t 75pw        sq ~�ήCUq ~ q ~�9t 1490t 84pw@5oz�G�sq ~�ήCtq ~ q ~�9t 1491t 75pw        sq ~�ήCq ~ q ~�9t 1491t 84pw@5oz�G�sq ~�ήC"�q ~ q ~�9t 1492t 84pw@5oz�G�sq ~�ήC&�q ~ q ~�9t 1493t 84pw@@�鹙�sq ~�ήC"zq ~ q ~�9t 1494t 61pw        sq ~�ήC*Yq ~ q ~�9t 1494t 84pw@5oz�G�sq ~�ήC.q ~ q ~�9t 1495t 84pw@5oz�G�sq ~�ήC.9q ~ q ~�9t 1496t 75pw        sq ~�ήC1�q ~ q ~�9t 1496t 84pw@#�k�(&sq ~�ήC-�q ~ q ~�9t 1497t 61pw        sq ~�ήC5�q ~ q ~�9t 1497t 84pw@@�鹙�sq ~�ήC9]q ~ q ~�9t 1498t 84pw@@�鹙�sq ~�ήC9|q ~ q ~�9t 1499t 75pw        sq ~�ήC=q ~ q ~�9t 1499t 84pw@$      sq ~��W�{�q ~ q ~�9t 15t 0pw        sq ~��W�3�q ~ q ~�9t 15t 12pw@8�H��fhsq ~��W�4vq ~ q ~�9t 15t 16pw@$      sq ~��W�7�q ~ q ~�9t 15t 22pw@3�~�]|sq ~��W�7�q ~ q ~�9t 15t 23pw@$sj�a'sq ~��W�|(q ~ q ~�9t 15t 3pw@ ,걉��sq ~��W�<q ~ q ~�9t 15t 37pw@$�(�>8sq ~��W�|�q ~ q ~�9t 15t 7pw��|#�]v�sq ~��Zy��q ~ q ~�9t 150t 84pw@$      sq ~�ήMq ~ q ~�9t 1500t 84pw@F�U�i�sq ~�ήMaq ~ q ~�9t 1501t 61pw        sq ~�ήM@q ~ q ~�9t 1501t 84pw@$      sq ~�ήM"q ~ q ~�9t 1502t 61pw        sq ~�ήM#q ~ q ~�9t 1502t 84pw@@�鹙�sq ~�ήM&�q ~ q ~�9t 1503t 84pw@5oz�G�sq ~�ήM"�q ~ q ~�9t 1504t 61pw        sq ~�ήM*�q ~ q ~�9t 1504t 84pw@5oz�G�sq ~�ήM&eq ~ q ~�9t 1505t 61pw        sq ~�ήM.Dq ~ q ~�9t 1505t 84pw@$      sq ~�ήM.cq ~ q ~�9t 1506t 75pw        sq ~�ήM2q ~ q ~�9t 1506t 84pw@5oz�G�sq ~�ήM-�q ~ q ~�9t 1507t 61pw        sq ~�ήM5�q ~ q ~�9t 1507t 84pw@$      sq ~�ήM5�q ~ q ~�9t 1508t 75pw        sq ~�ήM9�q ~ q ~�9t 1508t 84pw@@�鹙�sq ~�ήM9�q ~ q ~�9t 1509t 75pw        sq ~�ήM=Hq ~ q ~�9t 1509t 84pw@5oz�G�sq ~��Zy�q ~ q ~�9t 151t 75pw        sq ~��Zy��q ~ q ~�9t 151t 84pw@@�鹙�sq ~�ήM�<q ~ q ~�9t 1510t 75pw        sq ~�ήM��q ~ q ~�9t 1510t 84pw@5oz�G�sq ~�ήM��q ~ q ~�9t 1511t 75pw        sq ~�ήM��q ~ q ~�9t 1511t 84pw@@�鹙�sq ~�ήM��q ~ q ~�9t 1512t 75pw        sq ~�ήM�`q ~ q ~�9t 1512t 84pw@5oz�G�sq ~�ήM�!q ~ q ~�9t 1513t 84pw@5oz�G�sq ~�ήM�q ~ q ~�9t 1514t 61pw        sq ~�ήM��q ~ q ~�9t 1514t 84pw@5oz�G�sq ~�ήM�q ~ q ~�9t 1515t 75pw        sq ~�ήM��q ~ q ~�9t 1515t 84pw@$      sq ~�ήM��q ~ q ~�9t 1516t 75pw        sq ~�ήM�dq ~ q ~�9t 1516t 84pw@5oz�G�sq ~�ήM��q ~ q ~�9t 1517t 75pw        sq ~�ήM�%q ~ q ~�9t 1517t 84pw@$      sq ~�ήM�Dq ~ q ~�9t 1518t 75pw        sq ~�ήM��q ~ q ~�9t 1518t 84pw@@�鹙�sq ~�ήM��q ~ q ~�9t 1519t 61pw        sq ~�ήM��q ~ q ~�9t 1519t 84pw@5oz�G�sq ~��Zy��q ~ q ~�9t 152t 75pw        sq ~��Zy�iq ~ q ~�9t 152t 84pw@$      sq ~�ήN=q ~ q ~�9t 1520t 84pw@5oz�G�sq ~�ήN\q ~ q ~�9t 1521t 75pw        sq ~�ήN�q ~ q ~�9t 1521t 84pw@F�U�i�sq ~�ήN�q ~ q ~�9t 1522t 84pw@$      sq ~�ήN�q ~ q ~�9t 1523t 84pw@5oz�G�sq ~�ήNbq ~ q ~�9t 1524t 61pw        sq ~�ήNAq ~ q ~�9t 1524t 84pw@$      sq ~�ήN#q ~ q ~�9t 1525t 61pw        sq ~�ήNq ~ q ~�9t 1525t 84pw@F�U�i�sq ~�ήN�q ~ q ~�9t 1526t 61pw        sq ~�ήN�q ~ q ~�9t 1526t 84pw@5oz�G�sq ~�ήN�q ~ q ~�9t 1527t 61pw        sq ~�ήN�q ~ q ~�9t 1527t 84pw@@�鹙�sq ~�ήN"Eq ~ q ~�9t 1528t 84pw@@�鹙�sq ~�ήN&q ~ q ~�9t 1529t 84pw@$      sq ~��Zy�*q ~ q ~�9t 153t 84pw@5oz�G�sq ~�ήNp�q ~ q ~�9t 1530t 61pw        sq ~�ήNx�q ~ q ~�9t 1530t 84pw@$      sq ~�ήN|]q ~ q ~�9t 1531t 84pw@5oz�G�sq ~�ήN||q ~ q ~�9t 1532t 75pw        sq ~�ήN�q ~ q ~�9t 1532t 84pw@@�鹙�sq ~�ήN�=q ~ q ~�9t 1533t 75pw        sq ~�ήN��q ~ q ~�9t 1533t 84pw@5oz�G�sq ~�ήN��q ~ q ~�9t 1534t 84pw@5oz�G�sq ~�ήN��q ~ q ~�9t 1535t 61pw        sq ~�ήN�aq ~ q ~�9t 1535t 84pw@@�鹙�sq ~�ήN�"q ~ q ~�9t 1536t 84pw@5oz�G�sq ~�ήN��q ~ q ~�9t 1537t 84pw@5oz�G�sq ~�ήN��q ~ q ~�9t 1538t 84pw@$      sq ~�ήN��q ~ q ~�9t 1539t 75pw        sq ~�ήN�eq ~ q ~�9t 1539t 84pw@5oz�G�sq ~��Zy�Iq ~ q ~�9t 154t 75pw        sq ~��Zy��q ~ q ~�9t 154t 84pw@5oz�G�sq ~�ήN�Yq ~ q ~�9t 1540t 75pw        sq ~�ήN��q ~ q ~�9t 1540t 84pw@5oz�G�sq ~�ήN�q ~ q ~�9t 1541t 75pw        sq ~�ήN�q ~ q ~�9t 1541t 84pw@5oz�G�sq ~�ήN�}q ~ q ~�9t 1542t 84pw@@�鹙�sq ~�ήN�_q ~ q ~�9t 1543t 61pw        sq ~�ήN�>q ~ q ~�9t 1543t 84pw@@�鹙�sq ~�ήN�]q ~ q ~�9t 1544t 75pw        sq ~�ήN��q ~ q ~�9t 1544t 84pw@$      sq ~�ήN�q ~ q ~�9t 1545t 75pw        sq ~�ήN��q ~ q ~�9t 1545t 84pw@$      sq ~�ήN��q ~ q ~�9t 1546t 75pw        sq ~�ήO�q ~ q ~�9t 1546t 84pw@@�鹙�sq ~�ήN�cq ~ q ~�9t 1547t 61pw        sq ~�ήOBq ~ q ~�9t 1547t 84pw@6k����5sq ~�ήO$q ~ q ~�9t 1548t 61pw        sq ~�ήOq ~ q ~�9t 1548t 84pw@@�鹙�sq ~�ήO�q ~ q ~�9t 1549t 84pw@5oz�G�sq ~��Zy�
q ~ q ~�9t 155t 75pw        sq ~��Zy��q ~ q ~�9t 155t 84pw@5oz�G�sq ~�ήOY{q ~ q ~�9t 1550t 61pw        sq ~�ήOaZq ~ q ~�9t 1550t 84pw@5oz�G�sq ~�ήOayq ~ q ~�9t 1551t 75pw        sq ~�ήOeq ~ q ~�9t 1551t 84pw@$      sq ~�ήOh�q ~ q ~�9t 1552t 84pw@5oz�G�sq ~�ήOl�q ~ q ~�9t 1553t 84pw@@�鹙�sq ~�ήOl�q ~ q ~�9t 1554t 75pw        sq ~�ήOp^q ~ q ~�9t 1554t 84pw@5oz�G�sq ~�ήOp}q ~ q ~�9t 1555t 75pw        sq ~�ήOtq ~ q ~�9t 1555t 84pw@5oz�G�sq ~�ήOt>q ~ q ~�9t 1556t 75pw        sq ~�ήOw�q ~ q ~�9t 1556t 84pw@@�鹙�sq ~�ήO{�q ~ q ~�9t 1557t 84pw@5oz�G�sq ~�ήO{�q ~ q ~�9t 1558t 75pw        sq ~�ήObq ~ q ~�9t 1558t 84pw@@�鹙�sq ~�ήO�#q ~ q ~�9t 1559t 84pw@@�鹙�sq ~��Zy�mq ~ q ~�9t 156t 84pw@@�鹙�sq ~�ήOչq ~ q ~�9t 1560t 84pw@5oz�G�sq ~�ήO�zq ~ q ~�9t 1561t 84pw@5oz�G�sq ~�ήO�\q ~ q ~�9t 1562t 61pw        sq ~�ήO�;q ~ q ~�9t 1562t 84pw@$      sq ~�ήO��q ~ q ~�9t 1563t 84pw@@�鹙�sq ~�ήO�q ~ q ~�9t 1564t 84pw@5oz�G�sq ~�ήO��q ~ q ~�9t 1565t 75pw        sq ~�ήO�~q ~ q ~�9t 1565t 84pw@$      sq ~�ήO�?q ~ q ~�9t 1566t 84pw@$      sq ~�ήO�!q ~ q ~�9t 1567t 61pw        sq ~�ήO� q ~ q ~�9t 1567t 84pw@5oz�G�sq ~�ήO��q ~ q ~�9t 1568t 61pw        sq ~�ήO��q ~ q ~�9t 1568t 84pw@$      sq ~�ήO�q ~ q ~�9t 1569t 61pw        sq ~�ήO��q ~ q ~�9t 1569t 84pw@@�鹙�sq ~��Zy��q ~ q ~�9t 157t 75pw        sq ~��Zy�.q ~ q ~�9t 157t 84pw@F�U�i�sq ~�ήPFvq ~ q ~�9t 1570t 75pw        sq ~�ήPJq ~ q ~�9t 1570t 84pw@$      sq ~�ήPE�q ~ q ~�9t 1571t 61pw        sq ~�ήPM�q ~ q ~�9t 1571t 84pw@5oz�G�sq ~�ήPI�q ~ q ~�9t 1572t 61pw        sq ~�ήPQ�q ~ q ~�9t 1572t 84pw@5oz�G�sq ~�ήPQ�q ~ q ~�9t 1573t 75pw        sq ~�ήPU[q ~ q ~�9t 1573t 84pw@F�U�i�sq ~�ήPUzq ~ q ~�9t 1574t 75pw        sq ~�ήPYq ~ q ~�9t 1574t 84pw@@�鹙�sq ~�ήP\�q ~ q ~�9t 1575t 84pw@5oz�G�sq ~�ήP\�q ~ q ~�9t 1576t 75pw        sq ~�ήP`�q ~ q ~�9t 1576t 84pw@5oz�G�sq ~�ήP\�q ~ q ~�9t 1577t 61pw        sq ~�ήPd_q ~ q ~�9t 1577t 84pw@5oz�G�sq ~�ήPh q ~ q ~�9t 1578t 84pw@5oz�G�sq ~�ήPh?q ~ q ~�9t 1579t 75pw        sq ~�ήPk�q ~ q ~�9t 1579t 84pw@F�U�i�sq ~��Zy�q ~ q ~�9t 158t 61pw        sq ~��Zy��q ~ q ~�9t 158t 84pw@5oz�G�sq ~�ήP�wq ~ q ~�9t 1580t 84pw@$      sq ~�ήP�Yq ~ q ~�9t 1581t 61pw        sq ~�ήP�8q ~ q ~�9t 1581t 84pw@$      sq ~�ήP�Wq ~ q ~�9t 1582t 75pw        sq ~�ήP��q ~ q ~�9t 1582t 84pw@@�鹙�sq ~�ήP��q ~ q ~�9t 1583t 61pw        sq ~�ήPɺq ~ q ~�9t 1583t 84pw@5oz�G�sq ~�ήP�{q ~ q ~�9t 1584t 84pw@$      sq ~�ήP�]q ~ q ~�9t 1585t 61pw        sq ~�ήP�<q ~ q ~�9t 1585t 84pw@@�鹙�sq ~�ήP�q ~ q ~�9t 1586t 61pw        sq ~�ήP��q ~ q ~�9t 1586t 84pw@5oz�G�sq ~�ήP��q ~ q ~�9t 1587t 61pw        sq ~�ήPؾq ~ q ~�9t 1587t 84pw@@�鹙�sq ~�ήPԠq ~ q ~�9t 1588t 61pw        sq ~�ήP�q ~ q ~�9t 1588t 84pw@5oz�G�sq ~�ήP�@q ~ q ~�9t 1589t 84pw@@�鹙�sq ~��Zy�q ~ q ~�9t 159t 75pw        sq ~��Zy��q ~ q ~�9t 159t 84pw@@�鹙�sq ~�ήQ2�q ~ q ~�9t 1590t 84pw@F�U�i�sq ~�ήQ.�q ~ q ~�9t 1591t 61pw        sq ~�ήQ6�q ~ q ~�9t 1591t 84pw@5oz�G�sq ~�ήQ6�q ~ q ~�9t 1592t 75pw        sq ~�ήQ:Xq ~ q ~�9t 1592t 84pw@$      sq ~�ήQ:wq ~ q ~�9t 1593t 75pw        sq ~�ήQ>q ~ q ~�9t 1593t 84pw@5oz�G�sq ~�ήQ>8q ~ q ~�9t 1594t 75pw        sq ~�ήQA�q ~ q ~�9t 1594t 84pw@5oz�G�sq ~�ήQE�q ~ q ~�9t 1595t 84pw@@�鹙�sq ~�ήQA}q ~ q ~�9t 1596t 61pw        sq ~�ήQI\q ~ q ~�9t 1596t 84pw@5oz�G�sq ~�ήQI{q ~ q ~�9t 1597t 75pw        sq ~�ήQMq ~ q ~�9t 1597t 84pw@$      sq ~�ήQP�q ~ q ~�9t 1598t 84pw@@�鹙�sq ~�ήQT�q ~ q ~�9t 1599t 84pw@5oz�G�sq ~��W�8Vq ~ q ~�9t 16t 17pw        sq ~��W�Nq ~ q ~�9t 16t 70pw@@�鹙�sq ~��Zy��q ~ q ~�9t 160t 75pw        sq ~��ZzFq ~ q ~�9t 160t 84pw@@�鹙�sq ~�ή[3 q ~ q ~�9t 1600t 84pw@@�鹙�sq ~�ή[6�q ~ q ~�9t 1601t 84pw@$      sq ~�ή[:�q ~ q ~�9t 1602t 84pw@@�鹙�sq ~�ή[:�q ~ q ~�9t 1603t 75pw        sq ~�ή[>Cq ~ q ~�9t 1603t 84pw@5oz�G�sq ~�ή[>bq ~ q ~�9t 1604t 75pw        sq ~�ή[Bq ~ q ~�9t 1604t 84pw@5oz�G�sq ~�ή[B#q ~ q ~�9t 1605t 75pw        sq ~�ή[E�q ~ q ~�9t 1605t 84pw@$      sq ~�ή[E�q ~ q ~�9t 1606t 75pw        sq ~�ή[I�q ~ q ~�9t 1606t 84pw@5oz�G�sq ~�ή[MGq ~ q ~�9t 1607t 84pw@5oz�G�sq ~�ή[Qq ~ q ~�9t 1608t 84pw@5oz�G�sq ~�ή[T�q ~ q ~�9t 1609t 84pw@@�鹙�sq ~��Zzeq ~ q ~�9t 161t 75pw        sq ~��Zzq ~ q ~�9t 161t 84pw@@�鹙�sq ~�ή[�_q ~ q ~�9t 1610t 84pw@$      sq ~�ή[� q ~ q ~�9t 1611t 84pw@5oz�G�sq ~�ή[�q ~ q ~�9t 1612t 61pw        sq ~�ή[��q ~ q ~�9t 1612t 84pw@@�鹙�sq ~�ή[��q ~ q ~�9t 1613t 84pw@@�鹙�sq ~�ή[��q ~ q ~�9t 1614t 75pw        sq ~�ή[�cq ~ q ~�9t 1614t 84pw@5oz�G�sq ~�ή[�Eq ~ q ~�9t 1615t 61pw        sq ~�ή[�$q ~ q ~�9t 1615t 84pw@5oz�G�sq ~�ή[�q ~ q ~�9t 1616t 61pw        sq ~�ή[��q ~ q ~�9t 1616t 84pw@5oz�G�sq ~�ή[��q ~ q ~�9t 1617t 61pw        sq ~�ή[��q ~ q ~�9t 1617t 84pw@@�鹙�sq ~�ή[�gq ~ q ~�9t 1618t 84pw@@�鹙�sq ~�ή[ņq ~ q ~�9t 1619t 75pw        sq ~�ή[�(q ~ q ~�9t 1619t 84pw@$      sq ~��Zz&q ~ q ~�9t 162t 75pw        sq ~��Zz�q ~ q ~�9t 162t 84pw@5oz�G�sq ~�ή\�q ~ q ~�9t 1620t 61pw        sq ~�ή\�q ~ q ~�9t 1620t 84pw@F�U�i�sq ~�ή\�q ~ q ~�9t 1621t 75pw        sq ~�ή\q ~ q ~�9t 1621t 84pw@5oz�G�sq ~�ή\aq ~ q ~�9t 1622t 61pw        sq ~�ή\#@q ~ q ~�9t 1622t 84pw@@�鹙�sq ~�ή\#_q ~ q ~�9t 1623t 75pw        sq ~�ή\'q ~ q ~�9t 1623t 84pw@5oz�G�sq ~�ή\' q ~ q ~�9t 1624t 75pw        sq ~�ή\*�q ~ q ~�9t 1624t 84pw@@�鹙�sq ~�ή\*�q ~ q ~�9t 1625t 75pw        sq ~�ή\.�q ~ q ~�9t 1625t 84pw@5oz�G�sq ~�ή\*eq ~ q ~�9t 1626t 61pw        sq ~�ή\2Dq ~ q ~�9t 1626t 84pw@F�U�i�sq ~�ή\6q ~ q ~�9t 1627t 84pw@$      sq ~�ή\9�q ~ q ~�9t 1628t 84pw@5oz�G�sq ~�ή\9�q ~ q ~�9t 1629t 75pw        sq ~�ή\=�q ~ q ~�9t 1629t 84pw@$      sq ~��Zz�q ~ q ~�9t 163t 84pw@5oz�G�sq ~�ή\�{q ~ q ~�9t 1630t 75pw        sq ~�ή\�q ~ q ~�9t 1630t 84pw@@�鹙�sq ~�ή\��q ~ q ~�9t 1631t 84pw@5oz�G�sq ~�ή\��q ~ q ~�9t 1632t 61pw        sq ~�ή\��q ~ q ~�9t 1632t 84pw@@�鹙�sq ~�ή\�`q ~ q ~�9t 1633t 84pw@F�U�i�sq ~�ή\�q ~ q ~�9t 1634t 75pw        sq ~�ή\�!q ~ q ~�9t 1634t 84pw@$      sq ~�ή\�q ~ q ~�9t 1635t 61pw        sq ~�ή\��q ~ q ~�9t 1635t 84pw@@�鹙�sq ~�ή\��q ~ q ~�9t 1636t 61pw        sq ~�ή\��q ~ q ~�9t 1636t 84pw@@�鹙�sq ~�ή\�dq ~ q ~�9t 1637t 84pw@@�鹙�sq ~�ή\��q ~ q ~�9t 1638t 75pw        sq ~�ή\�%q ~ q ~�9t 1638t 84pw@$      sq ~�ή\�Dq ~ q ~�9t 1639t 75pw        sq ~�ή\��q ~ q ~�9t 1639t 84pw@$      sq ~��Zzkq ~ q ~�9t 164t 61pw        sq ~��ZzJq ~ q ~�9t 164t 84pw@$      sq ~�ή\��q ~ q ~�9t 1640t 61pw        sq ~�ή]|q ~ q ~�9t 1640t 84pw@$      sq ~�ή]�q ~ q ~�9t 1641t 75pw        sq ~�ή]=q ~ q ~�9t 1641t 84pw@5oz�G�sq ~�ή]�q ~ q ~�9t 1642t 84pw@@�鹙�sq ~�ή]�q ~ q ~�9t 1643t 61pw        sq ~�ή]�q ~ q ~�9t 1643t 84pw@@�鹙�sq ~�ή]�q ~ q ~�9t 1644t 75pw        sq ~�ή]�q ~ q ~�9t 1644t 84pw@F�U�i�sq ~�ή]Aq ~ q ~�9t 1645t 84pw@$      sq ~�ή]q ~ q ~�9t 1646t 84pw@5oz�G�sq ~�ή]!q ~ q ~�9t 1647t 75pw        sq ~�ή]�q ~ q ~�9t 1647t 84pw@5oz�G�sq ~�ή]"�q ~ q ~�9t 1648t 84pw@@�鹙�sq ~�ή]&Eq ~ q ~�9t 1649t 84pw@$      sq ~��Zz,q ~ q ~�9t 165t 61pw        sq ~��Zzq ~ q ~�9t 165t 84pw@F�U�i�sq ~�ή]p�q ~ q ~�9t 1650t 61pw        sq ~�ή]x�q ~ q ~�9t 1650t 84pw@@�鹙�sq ~�ή]t�q ~ q ~�9t 1651t 61pw        sq ~�ή]|�q ~ q ~�9t 1651t 84pw@5oz�G�sq ~�ή]�]q ~ q ~�9t 1652t 84pw@M]��%��sq ~�ή]�|q ~ q ~�9t 1653t 75pw        sq ~�ή]�q ~ q ~�9t 1653t 84pw@$      sq ~�ή]�=q ~ q ~�9t 1654t 75pw        sq ~�ή]��q ~ q ~�9t 1654t 84pw@5oz�G�sq ~�ή]��q ~ q ~�9t 1655t 75pw        sq ~�ή]��q ~ q ~�9t 1655t 84pw@5oz�G�sq ~�ή]�aq ~ q ~�9t 1656t 84pw@5oz�G�sq ~�ή]�"q ~ q ~�9t 1657t 84pw@@�鹙�sq ~�ή]��q ~ q ~�9t 1658t 84pw@5oz�G�sq ~�ή]��q ~ q ~�9t 1659t 61pw        sq ~�ή]��q ~ q ~�9t 1659t 84pw@M]��%��sq ~��Zz�q ~ q ~�9t 166t 61pw        sq ~��Zz�q ~ q ~�9t 166t 84pw@F�U�i�sq ~�ή]�q ~ q ~�9t 1660t 75pw        sq ~�ή]�:q ~ q ~�9t 1660t 84pw@@�鹙�sq ~�ή]�q ~ q ~�9t 1661t 61pw        sq ~�ή]��q ~ q ~�9t 1661t 84pw@5oz�G�sq ~�ή]��q ~ q ~�9t 1662t 84pw@$      sq ~�ή]�}q ~ q ~�9t 1663t 84pw@$      sq ~�ή]�>q ~ q ~�9t 1664t 84pw@&5�k�sq ~�ή]� q ~ q ~�9t 1665t 61pw        sq ~�ή]��q ~ q ~�9t 1665t 84pw@@�鹙�sq ~�ή^�q ~ q ~�9t 1666t 84pw@F�U�i�sq ~�ή]��q ~ q ~�9t 1667t 61pw        sq ~�ή^�q ~ q ~�9t 1667t 84pw@$      sq ~�ή^�q ~ q ~�9t 1668t 75pw        sq ~�ή^Bq ~ q ~�9t 1668t 84pw@5oz�G�sq ~�ή^q ~ q ~�9t 1669t 84pw@@�鹙�sq ~��Zz�q ~ q ~�9t 167t 75pw        sq ~��Zz�q ~ q ~�9t 167t 84pw@@�鹙�sq ~�ή^]�q ~ q ~�9t 1670t 75pw        sq ~�ή^a�q ~ q ~�9t 1670t 84pw@@�鹙�sq ~�ή^eZq ~ q ~�9t 1671t 84pw@F�U�i�sq ~�ή^eyq ~ q ~�9t 1672t 75pw        sq ~�ή^iq ~ q ~�9t 1672t 84pw@5oz�G�sq ~�ή^l�q ~ q ~�9t 1673t 84pw@5oz�G�sq ~�ή^l�q ~ q ~�9t 1674t 75pw        sq ~�ή^p�q ~ q ~�9t 1674t 84pw@$      sq ~�ή^lq ~ q ~�9t 1675t 61pw        sq ~�ή^t^q ~ q ~�9t 1675t 84pw@5oz�G�sq ~�ή^p@q ~ q ~�9t 1676t 61pw        sq ~�ή^xq ~ q ~�9t 1676t 84pw@5oz�G�sq ~�ή^{�q ~ q ~�9t 1677t 84pw@5oz�G�sq ~�ή^{�q ~ q ~�9t 1678t 75pw        sq ~�ή^�q ~ q ~�9t 1678t 84pw@5oz�G�sq ~�ή^�bq ~ q ~�9t 1679t 84pw@$      sq ~��Zz�q ~ q ~�9t 168t 75pw        sq ~��ZzNq ~ q ~�9t 168t 84pw@$      sq ~�ή^��q ~ q ~�9t 1680t 84pw@5oz�G�sq ~�ή^�q ~ q ~�9t 1681t 75pw        sq ~�ή^ٹq ~ q ~�9t 1681t 84pw@5oz�G�sq ~�ή^�zq ~ q ~�9t 1682t 84pw@$      sq ~�ή^�\q ~ q ~�9t 1683t 61pw        sq ~�ή^�;q ~ q ~�9t 1683t 84pw@5oz�G�sq ~�ή^��q ~ q ~�9t 1684t 84pw@F�U�i�sq ~�ή^�q ~ q ~�9t 1685t 84pw@@�鹙�sq ~�ή^�q ~ q ~�9t 1686t 61pw        sq ~�ή^�~q ~ q ~�9t 1686t 84pw@@�鹙�sq ~�ή^�?q ~ q ~�9t 1687t 84pw@$O,5/*�sq ~�ή^� q ~ q ~�9t 1688t 84pw@@�鹙�sq ~�ή^��q ~ q ~�9t 1689t 61pw        sq ~�ή^��q ~ q ~�9t 1689t 84pw@5oz�G�sq ~��Zzmq ~ q ~�9t 169t 75pw        sq ~��Zz#q ~ q ~�9t 169t 84pw@@�鹙�sq ~�ή_JWq ~ q ~�9t 1690t 84pw@5oz�G�sq ~�ή_Nq ~ q ~�9t 1691t 84pw@$      sq ~�ή_N7q ~ q ~�9t 1692t 75pw        sq ~�ή_Q�q ~ q ~�9t 1692t 84pw@@�鹙�sq ~�ή_M�q ~ q ~�9t 1693t 61pw        sq ~�ή_U�q ~ q ~�9t 1693t 84pw@F�U�i�sq ~�ή_Q|q ~ q ~�9t 1694t 61pw        sq ~�ή_Y[q ~ q ~�9t 1694t 84pw@@�鹙�sq ~�ή_]q ~ q ~�9t 1695t 84pw@$      sq ~�ή_X�q ~ q ~�9t 1696t 61pw        sq ~�ή_`�q ~ q ~�9t 1696t 84pw@5oz�G�sq ~�ή_d�q ~ q ~�9t 1697t 84pw@5oz�G�sq ~�ή_d�q ~ q ~�9t 1698t 75pw        sq ~�ή_h_q ~ q ~�9t 1698t 84pw@$      sq ~�ή_h~q ~ q ~�9t 1699t 75pw        sq ~�ή_l q ~ q ~�9t 1699t 84pw@$      sq ~��W�;|q ~ q ~�9t 17t 12pw����R�sq ~��W�<6q ~ q ~�9t 17t 18pw        sq ~��W�@q ~ q ~�9t 17t 29pw@&�.��'�sq ~��Wă�q ~ q ~�9t 17t 3pw����Ȝ sq ~��W�G;q ~ q ~�9t 17t 46pw@/����fsq ~��Zzrq ~ q ~�9t 170t 75pw        sq ~��Zzu�q ~ q ~�9t 170t 84pw@F�U�i�sq ~�ήiJ�q ~ q ~�9t 1700t 84pw@$      sq ~�ήiNBq ~ q ~�9t 1701t 84pw@5oz�G�sq ~�ήiRq ~ q ~�9t 1702t 84pw@$      sq ~�ήiR"q ~ q ~�9t 1703t 75pw        sq ~�ήiU�q ~ q ~�9t 1703t 84pw@@�鹙�sq ~�ήiY�q ~ q ~�9t 1704t 84pw@$      sq ~�ήiUgq ~ q ~�9t 1705t 61pw        sq ~�ήi]Fq ~ q ~�9t 1705t 84pw@5oz�G�sq ~�ήiY(q ~ q ~�9t 1706t 61pw        sq ~�ήiaq ~ q ~�9t 1706t 84pw@5oz�G�sq ~�ήia&q ~ q ~�9t 1707t 75pw        sq ~�ήid�q ~ q ~�9t 1707t 84pw@5oz�G�sq ~�ήid�q ~ q ~�9t 1708t 75pw        sq ~�ήih�q ~ q ~�9t 1708t 84pw@$      sq ~�ήidkq ~ q ~�9t 1709t 61pw        sq ~�ήilJq ~ q ~�9t 1709t 84pw@$      sq ~��Zzu�q ~ q ~�9t 171t 75pw        sq ~��Zzyfq ~ q ~�9t 171t 84pw@$      sq ~�ήi��q ~ q ~�9t 1710t 84pw@5oz�G�sq ~�ήi¡q ~ q ~�9t 1711t 84pw@@�鹙�sq ~�ήi��q ~ q ~�9t 1712t 61pw        sq ~�ήi�bq ~ q ~�9t 1712t 84pw@$      sq ~�ήi�#q ~ q ~�9t 1713t 84pw@5oz�G�sq ~�ήi�q ~ q ~�9t 1714t 61pw        sq ~�ήi��q ~ q ~�9t 1714t 84pw@$      sq ~�ήi��q ~ q ~�9t 1715t 61pw        sq ~�ήiѥq ~ q ~�9t 1715t 84pw@@�鹙�sq ~�ήi͇q ~ q ~�9t 1716t 61pw        sq ~�ήi�fq ~ q ~�9t 1716t 84pw@$      sq ~�ήi�'q ~ q ~�9t 1717t 84pw@$      sq ~�ήi��q ~ q ~�9t 1718t 84pw@F�U�i�sq ~�ήi�q ~ q ~�9t 1719t 84pw@F�U�i�sq ~��Zz}'q ~ q ~�9t 172t 84pw@5oz�G�sq ~�ήj/�q ~ q ~�9t 1720t 75pw        sq ~�ήj3?q ~ q ~�9t 1720t 84pw@F�U�i�sq ~�ήj/!q ~ q ~�9t 1721t 61pw        sq ~�ήj7 q ~ q ~�9t 1721t 84pw@5oz�G�sq ~�ήj:�q ~ q ~�9t 1722t 84pw@@�鹙�sq ~�ήj6�q ~ q ~�9t 1723t 61pw        sq ~�ήj>�q ~ q ~�9t 1723t 84pw@$      sq ~�ήj>�q ~ q ~�9t 1724t 75pw        sq ~�ήjBCq ~ q ~�9t 1724t 84pw@5oz�G�sq ~�ήjBbq ~ q ~�9t 1725t 75pw        sq ~�ήjFq ~ q ~�9t 1725t 84pw@"D�^���sq ~�ήjF#q ~ q ~�9t 1726t 75pw        sq ~�ήjI�q ~ q ~�9t 1726t 84pw@5oz�G�sq ~�ήjM�q ~ q ~�9t 1727t 84pw@@�鹙�sq ~�ήjIhq ~ q ~�9t 1728t 61pw        sq ~�ήjQGq ~ q ~�9t 1728t 84pw@$      sq ~�ήjM)q ~ q ~�9t 1729t 61pw        sq ~�ήjUq ~ q ~�9t 1729t 84pw@$      sq ~��Zz��q ~ q ~�9t 173t 84pw@@�鹙�sq ~�ήj��q ~ q ~�9t 1730t 75pw        sq ~�ήj��q ~ q ~�9t 1730t 84pw@$      sq ~�ήj��q ~ q ~�9t 1731t 61pw        sq ~�ήj�_q ~ q ~�9t 1731t 84pw@@�鹙�sq ~�ήj�Aq ~ q ~�9t 1732t 61pw        sq ~�ήj� q ~ q ~�9t 1732t 84pw@$      sq ~�ήj�q ~ q ~�9t 1733t 61pw        sq ~�ήj��q ~ q ~�9t 1733t 84pw@$      sq ~�ήj��q ~ q ~�9t 1734t 84pw@$      sq ~�ήj��q ~ q ~�9t 1735t 75pw        sq ~�ήj�cq ~ q ~�9t 1735t 84pw@@�鹙�sq ~�ήj��q ~ q ~�9t 1736t 75pw        sq ~�ήj�$q ~ q ~�9t 1736t 84pw@$      sq ~�ήj�q ~ q ~�9t 1737t 61pw        sq ~�ήj��q ~ q ~�9t 1737t 84pw@$      sq ~�ήj��q ~ q ~�9t 1738t 61pw        sq ~�ήjŦq ~ q ~�9t 1738t 84pw@$      sq ~�ήj��q ~ q ~�9t 1739t 61pw        sq ~�ήj�gq ~ q ~�9t 1739t 84pw@@�鹙�sq ~��Zz�q ~ q ~�9t 174t 75pw        sq ~��Zz��q ~ q ~�9t 174t 84pw@@�鹙�sq ~�ήk�q ~ q ~�9t 1740t 84pw@5oz�G�sq ~�ήk�q ~ q ~�9t 1741t 84pw@5oz�G�sq ~�ήk�q ~ q ~�9t 1742t 61pw        sq ~�ήk#q ~ q ~�9t 1742t 84pw@5oz�G�sq ~�ήkaq ~ q ~�9t 1743t 61pw        sq ~�ήk'@q ~ q ~�9t 1743t 84pw@5oz�G�sq ~�ήk#"q ~ q ~�9t 1744t 61pw        sq ~�ήk+q ~ q ~�9t 1744t 84pw@@�鹙�sq ~�ήk+ q ~ q ~�9t 1745t 75pw        sq ~�ήk.�q ~ q ~�9t 1745t 84pw@5y	=[ssq ~�ήk*�q ~ q ~�9t 1746t 61pw        sq ~�ήk2�q ~ q ~�9t 1746t 84pw@$      sq ~�ήk.eq ~ q ~�9t 1747t 61pw        sq ~�ήk6Dq ~ q ~�9t 1747t 84pw@5oz�G�sq ~�ήk:q ~ q ~�9t 1748t 84pw@5oz�G�sq ~�ήk=�q ~ q ~�9t 1749t 84pw@M]��%��sq ~��Zz��q ~ q ~�9t 175t 75pw        sq ~��Zz�jq ~ q ~�9t 175t 84pw@5oz�G�sq ~�ήk�}q ~ q ~�9t 1750t 61pw        sq ~�ήk�\q ~ q ~�9t 1750t 84pw@@�鹙�sq ~�ήk�>q ~ q ~�9t 1751t 61pw        sq ~�ήk�q ~ q ~�9t 1751t 84pw@5oz�G�sq ~�ήk�<q ~ q ~�9t 1752t 75pw        sq ~�ήk��q ~ q ~�9t 1752t 84pw@$      sq ~�ήk��q ~ q ~�9t 1753t 84pw@5oz�G�sq ~�ήk��q ~ q ~�9t 1754t 75pw        sq ~�ήk�`q ~ q ~�9t 1754t 84pw@@�鹙�sq ~�ήk�!q ~ q ~�9t 1755t 84pw@F�U�i�sq ~�ήk�@q ~ q ~�9t 1756t 75pw        sq ~�ήk��q ~ q ~�9t 1756t 84pw@$      sq ~�ήk��q ~ q ~�9t 1757t 84pw@5oz�G�sq ~�ήk��q ~ q ~�9t 1758t 61pw        sq ~�ήk�dq ~ q ~�9t 1758t 84pw@@�鹙�sq ~�ήk�%q ~ q ~�9t 1759t 84pw@$      sq ~��Zz��q ~ q ~�9t 176t 75pw        sq ~��Zz�+q ~ q ~�9t 176t 84pw@$      sq ~�ήlq ~ q ~�9t 1760t 75pw        sq ~�ήl�q ~ q ~�9t 1760t 84pw@5oz�G�sq ~�ήl|q ~ q ~�9t 1761t 84pw@@�鹙�sq ~�ήl=q ~ q ~�9t 1762t 84pw@5oz�G�sq ~�ήlq ~ q ~�9t 1763t 61pw        sq ~�ήl�q ~ q ~�9t 1763t 84pw@5oz�G�sq ~�ήlq ~ q ~�9t 1764t 75pw        sq ~�ήl�q ~ q ~�9t 1764t 84pw@$      sq ~�ήl�q ~ q ~�9t 1765t 75pw        sq ~�ήl�q ~ q ~�9t 1765t 84pw@@�鹙�sq ~�ήlAq ~ q ~�9t 1766t 84pw@@�鹙�sq ~�ήlq ~ q ~�9t 1767t 84pw@5oz�G�sq ~�ήl!q ~ q ~�9t 1768t 75pw        sq ~�ήl"�q ~ q ~�9t 1768t 84pw@5oz�G�sq ~�ήl�q ~ q ~�9t 1769t 61pw        sq ~�ήl&�q ~ q ~�9t 1769t 84pw@@�鹙�sq ~��Zz�q ~ q ~�9t 177t 61pw        sq ~��Zz��q ~ q ~�9t 177t 84pw@F�U�i�sq ~�ήlq;q ~ q ~�9t 1770t 61pw        sq ~�ήlyq ~ q ~�9t 1770t 84pw@$      sq ~�ήly9q ~ q ~�9t 1771t 75pw        sq ~�ήl|�q ~ q ~�9t 1771t 84pw@$      sq ~�ήlx�q ~ q ~�9t 1772t 61pw        sq ~�ήl��q ~ q ~�9t 1772t 84pw@@�鹙�sq ~�ήl|~q ~ q ~�9t 1773t 61pw        sq ~�ήl�]q ~ q ~�9t 1773t 84pw@5oz�G�sq ~�ήl�?q ~ q ~�9t 1774t 61pw        sq ~�ήl�q ~ q ~�9t 1774t 84pw@@�鹙�sq ~�ήl��q ~ q ~�9t 1775t 84pw@$      sq ~�ήl��q ~ q ~�9t 1776t 75pw        sq ~�ήl��q ~ q ~�9t 1776t 84pw@5oz�G�sq ~�ήl��q ~ q ~�9t 1777t 61pw        sq ~�ήl�aq ~ q ~�9t 1777t 84pw@@�鹙�sq ~�ήl�Cq ~ q ~�9t 1778t 61pw��l|�1��sq ~�ήl��q ~ q ~�9t 1778t 75pw        sq ~�ήl�"q ~ q ~�9t 1778t 84pw@"9�{�1�sq ~�ήl�Aq ~ q ~�9t 1779t 75pw        sq ~�ήl��q ~ q ~�9t 1779t 84pw@5oz�G�sq ~��Zz��q ~ q ~�9t 178t 84pw@5oz�G�sq ~�ήl�q ~ q ~�9t 1780t 61pw        sq ~�ήl�yq ~ q ~�9t 1780t 84pw@5oz�G�sq ~�ήl�:q ~ q ~�9t 1781t 84pw@$      sq ~�ήl�q ~ q ~�9t 1782t 61pw        sq ~�ήl��q ~ q ~�9t 1782t 84pw@$      sq ~�ήl��q ~ q ~�9t 1783t 84pw@@�鹙�sq ~�ήl�}q ~ q ~�9t 1784t 84pw@@�鹙�sq ~�ήm >q ~ q ~�9t 1785t 84pw@$      sq ~�ήl� q ~ q ~�9t 1786t 61pw        sq ~�ήm�q ~ q ~�9t 1786t 84pw@@�鹙�sq ~�ήl��q ~ q ~�9t 1787t 61pw        sq ~�ήm�q ~ q ~�9t 1787t 84pw@5oz�G�sq ~�ήm�q ~ q ~�9t 1788t 75pw        sq ~�ήm�q ~ q ~�9t 1788t 84pw@$      sq ~�ήmcq ~ q ~�9t 1789t 61pw        sq ~�ήmBq ~ q ~�9t 1789t 84pw@#y�Ƚsq ~��Zz�nq ~ q ~�9t 179t 84pw@5oz�G�sq ~�ήm^6q ~ q ~�9t 1790t 75pw        sq ~�ήma�q ~ q ~�9t 1790t 84pw@@�鹙�sq ~�ήme�q ~ q ~�9t 1791t 84pw@@�鹙�sq ~�ήme�q ~ q ~�9t 1792t 75pw        sq ~�ήmiZq ~ q ~�9t 1792t 84pw@@�鹙�sq ~�ήmiyq ~ q ~�9t 1793t 75pw        sq ~�ήmmq ~ q ~�9t 1793t 84pw@$      sq ~�ήmm:q ~ q ~�9t 1794t 75pw        sq ~�ήmp�q ~ q ~�9t 1794t 84pw@@�鹙�sq ~�ήml�q ~ q ~�9t 1795t 61pw        sq ~�ήmt�q ~ q ~�9t 1795t 84pw@$      sq ~�ήmpq ~ q ~�9t 1796t 61pw        sq ~�ήmx^q ~ q ~�9t 1796t 84pw@@�鹙�sq ~�ήm|q ~ q ~�9t 1797t 84pw@>�wV�Asq ~�ήm�q ~ q ~�9t 1798t 84pw@5oz�G�sq ~�ήm��q ~ q ~�9t 1799t 84pw@@�鹙�sq ~��W�@q ~ q ~�9t 18t 19pw@-~a��.asq ~��W�F�q ~ q ~�9t 18t 33pw����#��sq ~��W�R!q ~ q ~�9t 18t 63pw�xQ�=��sq ~��Zz�bq ~ q ~�9t 180t 75pw        sq ~��Zz�q ~ q ~�9t 180t 84pw@5oz�G�sq ~�ήwZ#q ~ q ~�9t 1800t 61pw        sq ~�ήwbq ~ q ~�9t 1800t 84pw@$      sq ~�ήwb!q ~ q ~�9t 1801t 75pw        sq ~�ήwe�q ~ q ~�9t 1801t 84pw@@�鹙�sq ~�ήwi�q ~ q ~�9t 1802t 84pw@5oz�G�sq ~�ήwmEq ~ q ~�9t 1803t 84pw@@�鹙�sq ~�ήwi'q ~ q ~�9t 1804t 61pw        sq ~�ήwqq ~ q ~�9t 1804t 84pw@F�U�i�sq ~�ήwq%q ~ q ~�9t 1805t 75pw        sq ~�ήwt�q ~ q ~�9t 1805t 84pw@$      sq ~�ήwx�q ~ q ~�9t 1806t 84pw@@�鹙�sq ~�ήwtjq ~ q ~�9t 1807t 61pw        sq ~�ήw|Iq ~ q ~�9t 1807t 84pw@$      sq ~�ήw�
q ~ q ~�9t 1808t 84pw@5oz�G�sq ~�ήw{�q ~ q ~�9t 1809t 61pw        sq ~�ήw��q ~ q ~�9t 1809t 84pw@$      sq ~��Zz��q ~ q ~�9t 181t 61pw        sq ~��Zz��q ~ q ~�9t 181t 84pw@5oz�G�sq ~�ήw΂q ~ q ~�9t 1810t 61pw        sq ~�ήw�aq ~ q ~�9t 1810t 84pw@5oz�G�sq ~�ήw�"q ~ q ~�9t 1811t 84pw@$      sq ~�ήw�Aq ~ q ~�9t 1812t 75pw        sq ~�ήw��q ~ q ~�9t 1812t 84pw@%�]�7�sq ~�ήw�q ~ q ~�9t 1813t 75pw        sq ~�ήw�q ~ q ~�9t 1813t 84pw@@�鹙�sq ~�ήw��q ~ q ~�9t 1814t 75pw        sq ~�ήw�eq ~ q ~�9t 1814t 84pw@$      sq ~�ήw�q ~ q ~�9t 1815t 75pw        sq ~�ήw�&q ~ q ~�9t 1815t 84pw@F�U�i�sq ~�ήw�Eq ~ q ~�9t 1816t 75pw        sq ~�ήw��q ~ q ~�9t 1816t 84pw@#�)6I�sq ~�ήw��q ~ q ~�9t 1817t 61pw        sq ~�ήw�q ~ q ~�9t 1817t 84pw@$      sq ~�ήw�iq ~ q ~�9t 1818t 84pw@5oz�G�sq ~�ήw�Kq ~ q ~�9t 1819t 61pw        sq ~�ήw�*q ~ q ~�9t 1819t 84pw@5oz�G�sq ~��Zz�q ~ q ~�9t 182t 61pw        sq ~��Zz�q ~ q ~�9t 182t 84pw@5oz�G�sq ~�ήxB�q ~ q ~�9t 1820t 61pw        sq ~�ήxJ�q ~ q ~�9t 1820t 84pw@5oz�G�sq ~�ήxJ�q ~ q ~�9t 1821t 75pw        sq ~�ήxN�q ~ q ~�9t 1821t 84pw@@�鹙�sq ~�ήxRBq ~ q ~�9t 1822t 84pw@5oz�G�sq ~�ήxRaq ~ q ~�9t 1823t 75pw        sq ~�ήxVq ~ q ~�9t 1823t 84pw@@�鹙�sq ~�ήxV"q ~ q ~�9t 1824t 75pw        sq ~�ήxY�q ~ q ~�9t 1824t 84pw@$      sq ~�ήx]�q ~ q ~�9t 1825t 84pw@5oz�G�sq ~�ήxaFq ~ q ~�9t 1826t 84pw@5oz�G�sq ~�ήxeq ~ q ~�9t 1827t 84pw@$      sq ~�ήxe&q ~ q ~�9t 1828t 75pw        sq ~�ήxh�q ~ q ~�9t 1828t 84pw@5oz�G�sq ~�ήxh�q ~ q ~�9t 1829t 75pw        sq ~�ήxl�q ~ q ~�9t 1829t 84pw@%�ذ�|
sq ~��Zz�hq ~ q ~�9t 183t 61pw        sq ~��Zz�Gq ~ q ~�9t 183t 84pw@5oz�G�sq ~�ήx�q ~ q ~�9t 1830t 84pw@$      sq ~�ήx�q ~ q ~�9t 1831t 61pw        sq ~�ήx��q ~ q ~�9t 1831t 84pw@5oz�G�sq ~�ήxơq ~ q ~�9t 1832t 84pw@F�U�i�sq ~�ήxq ~ q ~�9t 1833t 61pw        sq ~�ήx�bq ~ q ~�9t 1833t 84pw@5oz�G�sq ~�ήxʁq ~ q ~�9t 1834t 75pw        sq ~�ήx�#q ~ q ~�9t 1834t 84pw@5oz�G�sq ~�ήx��q ~ q ~�9t 1835t 84pw@$      sq ~�ήx��q ~ q ~�9t 1836t 61pw        sq ~�ήxեq ~ q ~�9t 1836t 84pw@@�鹙�sq ~�ήx��q ~ q ~�9t 1837t 75pw        sq ~�ήx�fq ~ q ~�9t 1837t 84pw@@�鹙�sq ~�ήx�'q ~ q ~�9t 1838t 84pw@@�鹙�sq ~�ήx�	q ~ q ~�9t 1839t 61pw        sq ~�ήx��q ~ q ~�9t 1839t 84pw@$      sq ~��Zz�q ~ q ~�9t 184t 84pw@F�U�i�sq ~�ήy3~q ~ q ~�9t 1840t 84pw@$      sq ~�ήy7?q ~ q ~�9t 1841t 84pw@5oz�G�sq ~�ήy7^q ~ q ~�9t 1842t 75pw        sq ~�ήy; q ~ q ~�9t 1842t 84pw@@�鹙�sq ~�ήy>�q ~ q ~�9t 1843t 84pw@$      sq ~�ήy>�q ~ q ~�9t 1844t 75pw        sq ~�ήyB�q ~ q ~�9t 1844t 84pw@$      sq ~�ήyFCq ~ q ~�9t 1845t 84pw@5oz�G�sq ~�ήyFbq ~ q ~�9t 1846t 75pw        sq ~�ήyJq ~ q ~�9t 1846t 84pw@5o8��sq ~�ήyE�q ~ q ~�9t 1847t 61pw        sq ~�ήyM�q ~ q ~�9t 1847t 84pw@$      sq ~�ήyM�q ~ q ~�9t 1848t 75pw        sq ~�ήyQ�q ~ q ~�9t 1848t 84pw@5oz�G�sq ~�ήyUGq ~ q ~�9t 1849t 84pw@F�U�i�sq ~��Zz�'q ~ q ~�9t 185t 75pw        sq ~��Zz��q ~ q ~�9t 185t 84pw@F�U�i�sq ~�ήy��q ~ q ~�9t 1850t 61pw        sq ~�ήy��q ~ q ~�9t 1850t 84pw@$      sq ~�ήy��q ~ q ~�9t 1851t 61pw        sq ~�ήy��q ~ q ~�9t 1851t 84pw@5oz�G�sq ~�ήy�_q ~ q ~�9t 1852t 84pw@5oz�G�sq ~�ήy� q ~ q ~�9t 1853t 84pw@5oz�G�sq ~�ήy�q ~ q ~�9t 1854t 61pw        sq ~�ήy��q ~ q ~�9t 1854t 84pw@F�U�i�sq ~�ήy��q ~ q ~�9t 1855t 84pw@M]��%��sq ~�ήy��q ~ q ~�9t 1856t 75pw        sq ~�ήy�cq ~ q ~�9t 1856t 84pw@5oz�G�sq ~�ήy�Eq ~ q ~�9t 1857t 61pw        sq ~�ήy�$q ~ q ~�9t 1857t 84pw@5oz�G�sq ~�ήy�Cq ~ q ~�9t 1858t 75pw        sq ~�ήy��q ~ q ~�9t 1858t 84pw@$      sq ~�ήyɦq ~ q ~�9t 1859t 84pw@@�鹙�sq ~��Zz��q ~ q ~�9t 186t 61pw        sq ~��Z{ �q ~ q ~�9t 186t 84pw@$      sq ~�ήz�q ~ q ~�9t 1860t 75pw        sq ~�ήz<q ~ q ~�9t 1860t 84pw@$      sq ~�ήz�q ~ q ~�9t 1861t 84pw@$      sq ~�ήz�q ~ q ~�9t 1862t 61pw        sq ~�ήz#�q ~ q ~�9t 1862t 84pw@@�鹙�sq ~�ήz�q ~ q ~�9t 1863t 61pw        sq ~�ήz'q ~ q ~�9t 1863t 84pw@$      sq ~�ήz+@q ~ q ~�9t 1864t 84pw@F�U�i�sq ~�ήz'"q ~ q ~�9t 1865t 61pw        sq ~�ήz/q ~ q ~�9t 1865t 84pw@@�鹙�sq ~�ήz2�q ~ q ~�9t 1866t 84pw@5oz�G�sq ~�ήz6�q ~ q ~�9t 1867t 84pw@$      sq ~�ήz:Dq ~ q ~�9t 1868t 84pw@$      sq ~�ήz>q ~ q ~�9t 1869t 84pw@@�鹙�sq ~��Z{ �q ~ q ~�9t 187t 75pw        sq ~��Z{Kq ~ q ~�9t 187t 84pw@F�U�i�sq ~�ήz��q ~ q ~�9t 1870t 75pw        sq ~�ήz��q ~ q ~�9t 1870t 84pw@5oz�G�sq ~�ήz�\q ~ q ~�9t 1871t 84pw@@�鹙�sq ~�ήz�q ~ q ~�9t 1872t 84pw@$      sq ~�ήz��q ~ q ~�9t 1873t 61pw        sq ~�ήz��q ~ q ~�9t 1873t 84pw@5oz�G�sq ~�ήz��q ~ q ~�9t 1874t 61pw        sq ~�ήz��q ~ q ~�9t 1874t 84pw@5oz�G�sq ~�ήz�`q ~ q ~�9t 1875t 84pw@@�鹙�sq ~�ήz�Bq ~ q ~�9t 1876t 61pw        sq ~�ήz�!q ~ q ~�9t 1876t 84pw@$      sq ~�ήz�q ~ q ~�9t 1877t 61pw        sq ~�ήz��q ~ q ~�9t 1877t 84pw@5oz�G�sq ~�ήz��q ~ q ~�9t 1878t 84pw@M]��%��sq ~�ήz�dq ~ q ~�9t 1879t 84pw@"D�^�v.sq ~��Z{ -q ~ q ~�9t 188t 61pw        sq ~��Z{q ~ q ~�9t 188t 84pw@@�鹙�sq ~�ή{�q ~ q ~�9t 1880t 84pw@$      sq ~�ή{ �q ~ q ~�9t 1881t 61pw        sq ~�ή{�q ~ q ~�9t 1881t 84pw@5oz�G�sq ~�ή{|q ~ q ~�9t 1882t 84pw@5oz�G�sq ~�ή{�q ~ q ~�9t 1883t 75pw        sq ~�ή{=q ~ q ~�9t 1883t 84pw@5oz�G�sq ~�ή{q ~ q ~�9t 1884t 61pw        sq ~�ή{�q ~ q ~�9t 1884t 84pw@5{�j}9sq ~�ή{�q ~ q ~�9t 1885t 61pw        sq ~�ή{�q ~ q ~�9t 1885t 84pw@$      sq ~�ή{�q ~ q ~�9t 1886t 84pw@@�鹙�sq ~�ή{bq ~ q ~�9t 1887t 61pw        sq ~�ή{Aq ~ q ~�9t 1887t 84pw@@�鹙�sq ~�ή{#q ~ q ~�9t 1888t 84pw@$      sq ~�ή{#!q ~ q ~�9t 1889t 75pw        sq ~�ή{&�q ~ q ~�9t 1889t 84pw@@�鹙�sq ~��Z{+q ~ q ~�9t 189t 75pw        sq ~��Z{�q ~ q ~�9t 189t 84pw@@�鹙�sq ~�ή{u�q ~ q ~�9t 1890t 75pw        sq ~�ή{yYq ~ q ~�9t 1890t 84pw@$      sq ~�ή{}q ~ q ~�9t 1891t 84pw@5oz�G�sq ~�ή{x�q ~ q ~�9t 1892t 61pw        sq ~�ή{��q ~ q ~�9t 1892t 84pw@@�鹙�sq ~�ή{|�q ~ q ~�9t 1893t 61pw        sq ~�ή{��q ~ q ~�9t 1893t 84pw@@�鹙�sq ~�ή{�~q ~ q ~�9t 1894t 61pw        sq ~�ή{�]q ~ q ~�9t 1894t 84pw@5oz�G�sq ~�ή{�q ~ q ~�9t 1895t 84pw@@�鹙�sq ~�ή{� q ~ q ~�9t 1896t 61pw        sq ~�ή{��q ~ q ~�9t 1896t 84pw@5oz�G�sq ~�ή{��q ~ q ~�9t 1897t 84pw@5oz�G�sq ~�ή{�aq ~ q ~�9t 1898t 84pw@@�鹙�sq ~�ή{��q ~ q ~�9t 1899t 75pw        sq ~�ή{�"q ~ q ~�9t 1899t 84pw@@�鹙�sq ~��W�F�q ~ q ~�9t 19t 20pw@@�鹙�sq ~��Z{^cq ~ q ~�9t 190t 84pw@@�鹙�sq ~�ή�q�q ~ q ~�9t 1900t 61pw        sq ~�ή�y�q ~ q ~�9t 1900t 84pw@@�鹙�sq ~�ή�y�q ~ q ~�9t 1901t 75pw        sq ~�ή�}Dq ~ q ~�9t 1901t 84pw@$      sq ~�ή�}cq ~ q ~�9t 1902t 75pw        sq ~�ή��q ~ q ~�9t 1902t 84pw@$      sq ~�ή���q ~ q ~�9t 1903t 84pw@5oz�G�sq ~�ή���q ~ q ~�9t 1904t 61pw        sq ~�ή���q ~ q ~�9t 1904t 84pw@$      sq ~�ή��Hq ~ q ~�9t 1905t 84pw@@�鹙�sq ~�ή��gq ~ q ~�9t 1906t 75pw        sq ~�ή��	q ~ q ~�9t 1906t 84pw@$      sq ~�ή��(q ~ q ~�9t 1907t 75pw        sq ~�ή���q ~ q ~�9t 1907t 84pw@$      sq ~�ή���q ~ q ~�9t 1908t 61pw        sq ~�ή���q ~ q ~�9t 1908t 84pw@$      sq ~�ή��mq ~ q ~�9t 1909t 61pw        sq ~�ή��Lq ~ q ~�9t 1909t 84pw@$      sq ~��Z{ZEq ~ q ~�9t 191t 61pw        sq ~��Z{b$q ~ q ~�9t 191t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1910t 61pw        sq ~�ή���q ~ q ~�9t 1910t 84pw@@�鹙�sq ~�ή���q ~ q ~�9t 1911t 61pw        sq ~�ή��q ~ q ~�9t 1911t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1912t 61pw        sq ~�ή��dq ~ q ~�9t 1912t 84pw@5oz�G�sq ~�ή��%q ~ q ~�9t 1913t 84pw@$      sq ~�ή��Dq ~ q ~�9t 1914t 75pw        sq ~�ή���q ~ q ~�9t 1914t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1915t 75pw        sq ~�ή� �q ~ q ~�9t 1915t 84pw@5oz�G�sq ~�ή�hq ~ q ~�9t 1916t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1917t 75pw        sq ~�ή�)q ~ q ~�9t 1917t 84pw@5oz�G�sq ~�ή�Hq ~ q ~�9t 1918t 75pw        sq ~�ή��q ~ q ~�9t 1918t 84pw@$      sq ~�ή�	q ~ q ~�9t 1919t 75pw        sq ~�ή��q ~ q ~�9t 1919t 84pw@5oz�G�sq ~��Z{^q ~ q ~�9t 192t 61pw        sq ~��Z{e�q ~ q ~�9t 192t 84pw@$      sq ~�ή�bAq ~ q ~�9t 1920t 84pw@5oz�G�sq ~�ή�fq ~ q ~�9t 1921t 84pw@5oz�G�sq ~�ή�i�q ~ q ~�9t 1922t 84pw@5oz�G�sq ~�ή�e�q ~ q ~�9t 1923t 61pw        sq ~�ή�m�q ~ q ~�9t 1923t 84pw@5oz�G�sq ~�ή�ifq ~ q ~�9t 1924t 61pw        sq ~�ή�qEq ~ q ~�9t 1924t 84pw@5oz�G�sq ~�ή�uq ~ q ~�9t 1925t 84pw@@�鹙�sq ~�ή�u%q ~ q ~�9t 1926t 75pw        sq ~�ή�x�q ~ q ~�9t 1926t 84pw@5oz�G�sq ~�ή�x�q ~ q ~�9t 1927t 75pw        sq ~�ή�|�q ~ q ~�9t 1927t 84pw@5oz�G�sq ~�ή��Iq ~ q ~�9t 1928t 84pw@$      sq ~�ή��hq ~ q ~�9t 1929t 75pw        sq ~�ή��
q ~ q ~�9t 1929t 84pw@@�鹙�sq ~��Z{fq ~ q ~�9t 193t 75pw        sq ~��Z{i�q ~ q ~�9t 193t 84pw@" ��C�sq ~�ή���q ~ q ~�9t 1930t 61pw        sq ~�ή�֠q ~ q ~�9t 1930t 84pw@$      sq ~�ή�ֿq ~ q ~�9t 1931t 75pw        sq ~�ή��aq ~ q ~�9t 1931t 84pw@@�鹙�sq ~�ή��Cq ~ q ~�9t 1932t 61pw        sq ~�ή��"q ~ q ~�9t 1932t 84pw@5oz�G�sq ~�ή���q ~ q ~�9t 1933t 84pw@$      sq ~�ή��q ~ q ~�9t 1934t 84pw@$      sq ~�ή��q ~ q ~�9t 1935t 61pw        sq ~�ή��eq ~ q ~�9t 1935t 84pw@5oz�G�sq ~�ή��&q ~ q ~�9t 1936t 84pw@@�鹙�sq ~�ή��Eq ~ q ~�9t 1937t 75pw        sq ~�ή���q ~ q ~�9t 1937t 84pw@#�pi[��sq ~�ή���q ~ q ~�9t 1938t 61pw        sq ~�ή���q ~ q ~�9t 1938t 84pw@F�U�i�sq ~�ή���q ~ q ~�9t 1939t 75pw        sq ~�ή��iq ~ q ~�9t 1939t 84pw@F�U�i�sq ~��Z{mgq ~ q ~�9t 194t 84pw@5oz�G�sq ~�ή�J�q ~ q ~�9t 1940t 84pw@F�U�i�sq ~�ή�F�q ~ q ~�9t 1941t 61pw        sq ~�ή�N�q ~ q ~�9t 1941t 84pw@5oz�G�sq ~�ή�N�q ~ q ~�9t 1942t 75pw        sq ~�ή�R�q ~ q ~�9t 1942t 84pw@5oz�G�sq ~�ή�VBq ~ q ~�9t 1943t 84pw@@�鹙�sq ~�ή�R$q ~ q ~�9t 1944t 61pw        sq ~�ή�Zq ~ q ~�9t 1944t 84pw@$      sq ~�ή�U�q ~ q ~�9t 1945t 61pw        sq ~�ή�]�q ~ q ~�9t 1945t 84pw@@�鹙�sq ~�ή�a�q ~ q ~�9t 1946t 84pw@$      sq ~�ή�]gq ~ q ~�9t 1947t 61pw        sq ~�ή�eFq ~ q ~�9t 1947t 84pw@5oz�G�sq ~�ή�a(q ~ q ~�9t 1948t 61pw        sq ~�ή�iq ~ q ~�9t 1948t 84pw@F�U�i�sq ~�ή�l�q ~ q ~�9t 1949t 84pw@@�鹙�sq ~��Z{m�q ~ q ~�9t 195t 75pw        sq ~��Z{q(q ~ q ~�9t 195t 84pw@$      sq ~�ή��q ~ q ~�9t 1950t 61pw        sq ~�ή��^q ~ q ~�9t 1950t 84pw@$      sq ~�ή��}q ~ q ~�9t 1951t 75pw        sq ~�ή��q ~ q ~�9t 1951t 84pw@F�U�i�sq ~�ή���q ~ q ~�9t 1952t 84pw@$      sq ~�ή�ʡq ~ q ~�9t 1953t 84pw@5oz�G�sq ~�ή��bq ~ q ~�9t 1954t 84pw@#��<U�+sq ~�ή��#q ~ q ~�9t 1955t 84pw@@�鹙�sq ~�ή���q ~ q ~�9t 1956t 84pw@$      sq ~�ή���q ~ q ~�9t 1957t 61pw        sq ~�ή�٥q ~ q ~�9t 1957t 84pw@5oz�G�sq ~�ή�Շq ~ q ~�9t 1958t 61pw        sq ~�ή��fq ~ q ~�9t 1958t 84pw@@�鹙�sq ~�ή�݅q ~ q ~�9t 1959t 75pw        sq ~�ή��'q ~ q ~�9t 1959t 84pw@5oz�G�sq ~��Z{qGq ~ q ~�9t 196t 75pw        sq ~��Z{t�q ~ q ~�9t 196t 84pw@$      sq ~�ή�0q ~ q ~�9t 1960t 75pw        sq ~�ή�3�q ~ q ~�9t 1960t 84pw@$      sq ~�ή�3�q ~ q ~�9t 1961t 75pw        sq ~�ή�7~q ~ q ~�9t 1961t 84pw@$      sq ~�ή�3`q ~ q ~�9t 1962t 61pw        sq ~�ή�;?q ~ q ~�9t 1962t 84pw@$      sq ~�ή�? q ~ q ~�9t 1963t 84pw@5oz�G�sq ~�ή�?q ~ q ~�9t 1964t 75pw        sq ~�ή�B�q ~ q ~�9t 1964t 84pw@5oz�G�sq ~�ή�F�q ~ q ~�9t 1965t 84pw@5oz�G�sq ~�ή�Bdq ~ q ~�9t 1966t 61pw        sq ~�ή�JCq ~ q ~�9t 1966t 84pw@@�鹙�sq ~�ή�Nq ~ q ~�9t 1967t 84pw@F�U�i�sq ~�ή�N#q ~ q ~�9t 1968t 75pw        sq ~�ή�Q�q ~ q ~�9t 1968t 84pw@@�鹙�sq ~�ή�U�q ~ q ~�9t 1969t 84pw@5oz�G�sq ~��Z{uq ~ q ~�9t 197t 75pw        sq ~��Z{x�q ~ q ~�9t 197t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1970t 84pw@5oz�G�sq ~�ή���q ~ q ~�9t 1971t 61pw        sq ~�ή���q ~ q ~�9t 1971t 84pw@5oz�G�sq ~�ή���q ~ q ~�9t 1972t 84pw@@�鹙�sq ~�ή���q ~ q ~�9t 1973t 61pw        sq ~�ή��_q ~ q ~�9t 1973t 84pw@5oz�G�sq ~�ή��Aq ~ q ~�9t 1974t 61pw        sq ~�ή�� q ~ q ~�9t 1974t 84pw@$      sq ~�ή��?q ~ q ~�9t 1975t 75pw        sq ~�ή���q ~ q ~�9t 1975t 84pw@$      sq ~�ή�� q ~ q ~�9t 1976t 75pw        sq ~�ή���q ~ q ~�9t 1976t 84pw@5oz�G�sq ~�ή��cq ~ q ~�9t 1977t 84pw@$��3�sq ~�ή�q ~ q ~�9t 1978t 75pw        sq ~�ή��$q ~ q ~�9t 1978t 84pw@5oz�G�sq ~�ή��Cq ~ q ~�9t 1979t 75pw        sq ~�ή���q ~ q ~�9t 1979t 84pw@$      sq ~��Z{x�q ~ q ~�9t 198t 75pw        sq ~��Z{|kq ~ q ~�9t 198t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1980t 61pw        sq ~�ή�{q ~ q ~�9t 1980t 84pw@$      sq ~�ή��q ~ q ~�9t 1981t 75pw        sq ~�ή� <q ~ q ~�9t 1981t 84pw@5oz�G�sq ~�ή�#�q ~ q ~�9t 1982t 84pw@@�鹙�sq ~�ή��q ~ q ~�9t 1983t 61pw        sq ~�ή�'�q ~ q ~�9t 1983t 84pw@5oz�G�sq ~�ή�'�q ~ q ~�9t 1984t 75pw        sq ~�ή�+q ~ q ~�9t 1984t 84pw@$      sq ~�ή�'aq ~ q ~�9t 1985t 61pw        sq ~�ή�/@q ~ q ~�9t 1985t 84pw@5oz�G�sq ~�ή�/_q ~ q ~�9t 1986t 75pw        sq ~�ή�3q ~ q ~�9t 1986t 84pw@5oz�G�sq ~�ή�3 q ~ q ~�9t 1987t 75pw        sq ~�ή�6�q ~ q ~�9t 1987t 84pw@5oz�G�sq ~�ή�:�q ~ q ~�9t 1988t 84pw@$      sq ~�ή�:�q ~ q ~�9t 1989t 75pw        sq ~�ή�>Dq ~ q ~�9t 1989t 84pw@@�鹙�sq ~��Z{�,q ~ q ~�9t 199t 84pw@5oz�G�sq ~�ή���q ~ q ~�9t 1990t 84pw@$      sq ~�ή���q ~ q ~�9t 1991t 61pw        sq ~�ή���q ~ q ~�9t 1991t 84pw@;4(�6�sq ~�ή��\q ~ q ~�9t 1992t 84pw@5oz�G�sq ~�ή��>q ~ q ~�9t 1993t 61pw        sq ~�ή��q ~ q ~�9t 1993t 84pw@F�U�i�sq ~�ή��<q ~ q ~�9t 1994t 75pw        sq ~�ή���q ~ q ~�9t 1994t 84pw@@�鹙�sq ~�ή���q ~ q ~�9t 1995t 84pw@$      sq ~�ή��`q ~ q ~�9t 1996t 84pw@@�鹙�sq ~�ή��!q ~ q ~�9t 1997t 84pw@$      sq ~�ή��@q ~ q ~�9t 1998t 75pw        sq ~�ή���q ~ q ~�9t 1998t 84pw@5oz�G�sq ~�ή��q ~ q ~�9t 1999t 75pw        sq ~�ή���q ~ q ~�9t 1999t 84pw@@�鹙�sq ~��W�*�q ~ q ~�9t 2t 2pw        sq ~��W�*�q ~ q ~�9t 2t 4pw@5oz�G�sq ~��W��eq ~ q ~�9t 2t 59pw@5oz�G�sq ~��Wř6q ~ q ~�9t 20t 21pw@*���{sq ~��Wř�q ~ q ~�9t 20t 26pw@(sj��bsq ~��W���q ~ q ~�9t 20t 4pw�k���9 sq ~��WŠ�q ~ q ~�9t 20t 42pw@$      sq ~��Wšq ~ q ~�9t 20t 44pw@'���#�sq ~��Z�Z�q ~ q ~�9t 200t 75pw        sq ~��Z�^�q ~ q ~�9t 200t 84pw@$      sq ~�ί�~�q ~ q ~�9t 2000t 84pw@5oz�G�sq ~�ί�z{q ~ q ~�9t 2001t 61pw        sq ~�ί��Zq ~ q ~�9t 2001t 84pw@5oz�G�sq ~�ί��yq ~ q ~�9t 2002t 75pw        sq ~�ί��q ~ q ~�9t 2002t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2003t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2004t 75pw        sq ~�ί���q ~ q ~�9t 2004t 84pw@$      sq ~�ί��q ~ q ~�9t 2005t 61pw        sq ~�ί��^q ~ q ~�9t 2005t 84pw@5oz�G�sq ~�ί��}q ~ q ~�9t 2006t 75pw        sq ~�ί��q ~ q ~�9t 2006t 84pw@5oz�G�sq ~�ί��>q ~ q ~�9t 2007t 75pw        sq ~�ί���q ~ q ~�9t 2007t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2008t 75pw        sq ~�ί���q ~ q ~�9t 2008t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2009t 61pw        sq ~�ί��bq ~ q ~�9t 2009t 84pw@F�U�i�sq ~��Z�bNq ~ q ~�9t 201t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2010t 84pw@$      sq ~�ί���q ~ q ~�9t 2011t 61pw        sq ~�ί���q ~ q ~�9t 2011t 84pw@5oz�G�sq ~�ί��zq ~ q ~�9t 2012t 84pw@$      sq ~�ί���q ~ q ~�9t 2013t 75pw        sq ~�ί��;q ~ q ~�9t 2013t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2014t 84pw@5oz�G�sq ~�ί�q ~ q ~�9t 2015t 75pw        sq ~�ί��q ~ q ~�9t 2015t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2016t 75pw        sq ~�ί�	~q ~ q ~�9t 2016t 84pw@5oz�G�sq ~�ί�	�q ~ q ~�9t 2017t 75pw        sq ~�ί�?q ~ q ~�9t 2017t 84pw@5oz�G�sq ~�ί�	!q ~ q ~�9t 2018t 61pw        sq ~�ί� q ~ q ~�9t 2018t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2019t 84pw@Q�"Ѱsq ~��Z�bmq ~ q ~�9t 202t 75pw        sq ~��Z�fq ~ q ~�9t 202t 84pw@F�U�i�sq ~�ί�_xq ~ q ~�9t 2020t 61pw        sq ~�ί�gWq ~ q ~�9t 2020t 84pw@@�鹙�sq ~�ί�c9q ~ q ~�9t 2021t 61pw        sq ~�ί�kq ~ q ~�9t 2021t 84pw@@�鹙�sq ~�ί�f�q ~ q ~�9t 2022t 61pw        sq ~�ί�n�q ~ q ~�9t 2022t 84pw@@�鹙�sq ~�ί�r�q ~ q ~�9t 2023t 84pw@$      sq ~�ί�n|q ~ q ~�9t 2024t 61pw        sq ~�ί�v[q ~ q ~�9t 2024t 84pw@@�鹙�sq ~�ί�vzq ~ q ~�9t 2025t 75pw        sq ~�ί�zq ~ q ~�9t 2025t 84pw@@�鹙�sq ~�ί�z;q ~ q ~�9t 2026t 75pw        sq ~�ί�}�q ~ q ~�9t 2026t 84pw@@�鹙�sq ~�ί�y�q ~ q ~�9t 2027t 61pw        sq ~�ί���q ~ q ~�9t 2027t 84pw@$      sq ~�ί���q ~ q ~�9t 2028t 75pw        sq ~�ί��_q ~ q ~�9t 2028t 84pw@$      sq ~�ί��Aq ~ q ~�9t 2029t 61pw        sq ~�ί�� q ~ q ~�9t 2029t 84pw@@�鹙�sq ~��Z�f.q ~ q ~�9t 203t 75pw        sq ~��Z�i�q ~ q ~�9t 203t 84pw@M]��%��sq ~�ί���q ~ q ~�9t 2030t 61pw        sq ~�ί�۶q ~ q ~�9t 2030t 84pw@$      sq ~�ί��wq ~ q ~�9t 2031t 84pw@5oz�G�sq ~�ί��8q ~ q ~�9t 2032t 84pw@@�鹙�sq ~�ί��Wq ~ q ~�9t 2033t 75pw        sq ~�ί���q ~ q ~�9t 2033t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2034t 75pw        sq ~�ί��q ~ q ~�9t 2034t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2035t 61pw        sq ~�ί��{q ~ q ~�9t 2035t 84pw@F�U�i�sq ~�ί��]q ~ q ~�9t 2036t 61pw        sq ~�ί��<q ~ q ~�9t 2036t 84pw@$      sq ~�ί��[q ~ q ~�9t 2037t 75pw        sq ~�ί���q ~ q ~�9t 2037t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2038t 75pw        sq ~�ί���q ~ q ~�9t 2038t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2039t 61pw        sq ~�ί��q ~ q ~�9t 2039t 84pw@$      sq ~��Z�m�q ~ q ~�9t 204t 84pw@5oz�G�sq ~�ί�Lsq ~ q ~�9t 2040t 75pw        sq ~�ί�Pq ~ q ~�9t 2040t 84pw@5oz�G�sq ~�ί�S�q ~ q ~�9t 2041t 84pw@5oz�G�sq ~�ί�O�q ~ q ~�9t 2042t 61pw        sq ~�ί�W�q ~ q ~�9t 2042t 84pw@@�鹙�sq ~�ί�Syq ~ q ~�9t 2043t 61pw        sq ~�ί�[Xq ~ q ~�9t 2043t 84pw@5oz�G�sq ~�ί�_q ~ q ~�9t 2044t 84pw@F�U�i�sq ~�ί�b�q ~ q ~�9t 2045t 84pw@@�鹙�sq ~�ί�^�q ~ q ~�9t 2046t 61pw        sq ~�ί�f�q ~ q ~�9t 2046t 84pw@@�鹙�sq ~�ί�f�q ~ q ~�9t 2047t 75pw        sq ~�ί�j\q ~ q ~�9t 2047t 84pw@5oz�G�sq ~�ί�j{q ~ q ~�9t 2048t 75pw        sq ~�ί�nq ~ q ~�9t 2048t 84pw@@�鹙�sq ~�ί�q�q ~ q ~�9t 2049t 84pw@5oz�G�sq ~��Z�qRq ~ q ~�9t 205t 84pw@$      sq ~�ί���q ~ q ~�9t 2050t 75pw        sq ~�ί��tq ~ q ~�9t 2050t 84pw@@�鹙�sq ~�ί�ēq ~ q ~�9t 2051t 75pw        sq ~�ί��5q ~ q ~�9t 2051t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2052t 61pw        sq ~�ί���q ~ q ~�9t 2052t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2053t 61pw        sq ~�ί�Ϸq ~ q ~�9t 2053t 84pw@$      sq ~�ί��xq ~ q ~�9t 2054t 84pw@5oz�G�sq ~�ί��Zq ~ q ~�9t 2055t 61pw        sq ~�ί��9q ~ q ~�9t 2055t 84pw@5oz�G�sq ~�ί��Xq ~ q ~�9t 2056t 75pw        sq ~�ί���q ~ q ~�9t 2056t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2057t 61pw        sq ~�ί�޻q ~ q ~�9t 2057t 84pw@5oz�G�sq ~�ί�ڝq ~ q ~�9t 2058t 61pw        sq ~�ί��|q ~ q ~�9t 2058t 84pw@$      sq ~�ί��^q ~ q ~�9t 2059t 61pw        sq ~�ί��=q ~ q ~�9t 2059t 84pw@$      sq ~��Z�qqq ~ q ~�9t 206t 75pw        sq ~��Z�uq ~ q ~�9t 206t 84pw@$      sq ~�ί�0�q ~ q ~�9t 2060t 61pw        sq ~�ί�8�q ~ q ~�9t 2060t 84pw@5oz�G�sq ~�ί�8�q ~ q ~�9t 2061t 75pw        sq ~�ί�<�q ~ q ~�9t 2061t 84pw@5oz�G�sq ~�ί�8vq ~ q ~�9t 2062t 61pw        sq ~�ί�@Uq ~ q ~�9t 2062t 84pw@5oz�G�sq ~�ί�Dq ~ q ~�9t 2063t 84pw@5oz�G�sq ~�ί�D5q ~ q ~�9t 2064t 75pw        sq ~�ί�G�q ~ q ~�9t 2064t 84pw@@�鹙�sq ~�ί�K�q ~ q ~�9t 2065t 84pw@F�U�i�sq ~�ί�Gzq ~ q ~�9t 2066t 61pw        sq ~�ί�OYq ~ q ~�9t 2066t 84pw@5oz�G�sq ~�ί�K;q ~ q ~�9t 2067t 61pw        sq ~�ί�Sq ~ q ~�9t 2067t 84pw@$      sq ~�ί�S9q ~ q ~�9t 2068t 75pw        sq ~�ί�V�q ~ q ~�9t 2068t 84pw@5oz�G�sq ~�ί�R�q ~ q ~�9t 2069t 61pw        sq ~�ί�Z�q ~ q ~�9t 2069t 84pw@%_?Jӕsq ~��Z�p�q ~ q ~�9t 207t 61pw        sq ~��Z�x�q ~ q ~�9t 207t 84pw@@�鹙�sq ~�ί��Sq ~ q ~�9t 2070t 61pw        sq ~�ί��2q ~ q ~�9t 2070t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2071t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2072t 75pw        sq ~�ί���q ~ q ~�9t 2072t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2073t 75pw        sq ~�ί��uq ~ q ~�9t 2073t 84pw@5oz�G�sq ~�ί��6q ~ q ~�9t 2074t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2075t 61pw        sq ~�ί���q ~ q ~�9t 2075t 84pw@F�U�i�sq ~�ί�øq ~ q ~�9t 2076t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2077t 75pw        sq ~�ί��yq ~ q ~�9t 2077t 84pw@5oz�G�sq ~�ί��:q ~ q ~�9t 2078t 84pw@5oz�G�sq ~�ί��Yq ~ q ~�9t 2079t 75pw        sq ~�ί���q ~ q ~�9t 2079t 84pw@5oz�G�sq ~��Z�x�q ~ q ~�9t 208t 75pw        sq ~��Z�|�q ~ q ~�9t 208t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2080t 61pw        sq ~�ί�!�q ~ q ~�9t 2080t 84pw@5oz�G�sq ~�ί�sq ~ q ~�9t 2081t 61pw        sq ~�ί�%Rq ~ q ~�9t 2081t 84pw@5oz�G�sq ~�ί�)q ~ q ~�9t 2082t 84pw@@�鹙�sq ~�ί�$�q ~ q ~�9t 2083t 61pw        sq ~�ί�,�q ~ q ~�9t 2083t 84pw@5oz�G�sq ~�ί�,�q ~ q ~�9t 2084t 75pw        sq ~�ί�0�q ~ q ~�9t 2084t 84pw@$      sq ~�ί�0�q ~ q ~�9t 2085t 75pw        sq ~�ί�4Vq ~ q ~�9t 2085t 84pw@5oz�G�sq ~�ί�8q ~ q ~�9t 2086t 84pw@$      sq ~�ί�86q ~ q ~�9t 2087t 75pw        sq ~�ί�;�q ~ q ~�9t 2087t 84pw@@�鹙�sq ~�ί�?�q ~ q ~�9t 2088t 84pw@5oz�G�sq ~�ί�CZq ~ q ~�9t 2089t 84pw@5oz�G�sq ~��Z�|�q ~ q ~�9t 209t 75pw        sq ~��Z��Vq ~ q ~�9t 209t 84pw@$      sq ~�ί��q ~ q ~�9t 2090t 61pw        sq ~�ί���q ~ q ~�9t 2090t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2091t 84pw@5oz�G�sq ~�ί��rq ~ q ~�9t 2092t 84pw@M]��%��sq ~�ί��3q ~ q ~�9t 2093t 84pw@$      sq ~�ί���q ~ q ~�9t 2094t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2095t 84pw@@�鹙�sq ~�ί��vq ~ q ~�9t 2096t 84pw@5oz�G�sq ~�ί��Xq ~ q ~�9t 2097t 61pw        sq ~�ί��7q ~ q ~�9t 2097t 84pw@%��_sq ~�ί��Vq ~ q ~�9t 2098t 75pw        sq ~�ί���q ~ q ~�9t 2098t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2099t 61pw        sq ~�ί���q ~ q ~�9t 2099t 84pw@5oz�G�sq ~��Wš�q ~ q ~�9t 21t 38pw@5oz�G�sq ~��Wťq ~ q ~�9t 21t 46pw        sq ~��Wť3q ~ q ~�9t 21t 47pw        sq ~��W���q ~ q ~�9t 21t 6pw        sq ~��Z���q ~ q ~�9t 210t 84pw@$      sq ~�ίɒxq ~ q ~�9t 2100t 75pw        sq ~�ίɖq ~ q ~�9t 2100t 84pw@F�U�i�sq ~�ίə�q ~ q ~�9t 2101t 84pw@@�鹙�sq ~�ίɕ�q ~ q ~�9t 2102t 61pw        sq ~�ίɝ�q ~ q ~�9t 2102t 84pw@5oz�G�sq ~�ίɡ]q ~ q ~�9t 2103t 84pw@5oz�G�sq ~�ίɡ|q ~ q ~�9t 2104t 75pw        sq ~�ίɥq ~ q ~�9t 2104t 84pw@5oz�G�sq ~�ίɨ�q ~ q ~�9t 2105t 84pw@5oz�G�sq ~�ίɤ�q ~ q ~�9t 2106t 61pw        sq ~�ίɬ�q ~ q ~�9t 2106t 84pw@$      sq ~�ίɰaq ~ q ~�9t 2107t 84pw@@�鹙�sq ~�ίɴ"q ~ q ~�9t 2108t 84pw@5oz�G�sq ~�ίɴAq ~ q ~�9t 2109t 75pw        sq ~�ίɷ�q ~ q ~�9t 2109t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 211t 61pw        sq ~��Z�֭q ~ q ~�9t 211t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2110t 75pw        sq ~�ί�
yq ~ q ~�9t 2110t 84pw@$      sq ~�ί�[q ~ q ~�9t 2111t 61pw        sq ~�ί�:q ~ q ~�9t 2111t 84pw@F�U�i�sq ~�ί�
q ~ q ~�9t 2112t 61pw        sq ~�ί��q ~ q ~�9t 2112t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2113t 61pw        sq ~�ί��q ~ q ~�9t 2113t 84pw@$      sq ~�ί�}q ~ q ~�9t 2114t 84pw@@�鹙�sq ~�ί�>q ~ q ~�9t 2115t 84pw@@�鹙�sq ~�ί� q ~ q ~�9t 2116t 61pw        sq ~�ί� �q ~ q ~�9t 2116t 84pw@5oz�G�sq ~�ί�!q ~ q ~�9t 2117t 75pw        sq ~�ί�$�q ~ q ~�9t 2117t 84pw@F�U�i�sq ~�ί�$�q ~ q ~�9t 2118t 75pw        sq ~�ί�(�q ~ q ~�9t 2118t 84pw@5oz�G�sq ~�ί�,Bq ~ q ~�9t 2119t 84pw@@�鹙�sq ~��Z�ҏq ~ q ~�9t 212t 61pw��:����.sq ~��Z��nq ~ q ~�9t 212t 84pw@��Ұ�
sq ~�ί�{6q ~ q ~�9t 2120t 75pw        sq ~�ί�~�q ~ q ~�9t 2120t 84pw@$      sq ~�ίʂ�q ~ q ~�9t 2121t 84pw@5oz�G�sq ~�ίʆZq ~ q ~�9t 2122t 84pw@$      sq ~�ίʂ<q ~ q ~�9t 2123t 61pw        sq ~�ίʊq ~ q ~�9t 2123t 84pw@@�鹙�sq ~�ίʍ�q ~ q ~�9t 2124t 84pw@5oz�G�sq ~�ίʑ�q ~ q ~�9t 2125t 84pw@5oz�G�sq ~�ίʕ^q ~ q ~�9t 2126t 84pw@%�e�_csq ~�ίʑ@q ~ q ~�9t 2127t 61pw        sq ~�ίʙq ~ q ~�9t 2127t 84pw@@�鹙�sq ~�ίʕq ~ q ~�9t 2128t 61pw        sq ~�ίʜ�q ~ q ~�9t 2128t 84pw@5oz�G�sq ~�ίʘ�q ~ q ~�9t 2129t 61pw        sq ~�ίʠ�q ~ q ~�9t 2129t 84pw@5oz�G�sq ~��Z��Pq ~ q ~�9t 213t 61pw        sq ~��Z��/q ~ q ~�9t 213t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2130t 75pw        sq ~�ί��7q ~ q ~�9t 2130t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2131t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2132t 61pw        sq ~�ί���q ~ q ~�9t 2132t 84pw@#�c�E'sq ~�ί���q ~ q ~�9t 2133t 75pw        sq ~�ί��zq ~ q ~�9t 2133t 84pw@$      sq ~�ί���q ~ q ~�9t 2134t 75pw        sq ~�ί�;q ~ q ~�9t 2134t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2135t 84pw@5oz�G�sq ~�ί�q ~ q ~�9t 2136t 75pw        sq ~�ί�	�q ~ q ~�9t 2136t 84pw@5oz�G�sq ~�ί�	�q ~ q ~�9t 2137t 75pw        sq ~�ί�~q ~ q ~�9t 2137t 84pw@$      sq ~�ί�?q ~ q ~�9t 2138t 84pw@5oz�G�sq ~�ί� q ~ q ~�9t 2139t 84pw@@�鹙�sq ~��Z��Nq ~ q ~�9t 214t 75pw        sq ~��Z���q ~ q ~�9t 214t 84pw@$      sq ~�ί�c�q ~ q ~�9t 2140t 75pw        sq ~�ί�g�q ~ q ~�9t 2140t 84pw@@�鹙�sq ~�ί�kWq ~ q ~�9t 2141t 84pw@F�U�i�sq ~�ί�g9q ~ q ~�9t 2142t 61pw        sq ~�ί�oq ~ q ~�9t 2142t 84pw@F�U�i�sq ~�ί�j�q ~ q ~�9t 2143t 61pw��l|�1�zsq ~�ί�r�q ~ q ~�9t 2143t 84pw@"9�{�1�sq ~�ί�r�q ~ q ~�9t 2144t 75pw        sq ~�ί�v�q ~ q ~�9t 2144t 84pw@5oz�G�sq ~�ί�v�q ~ q ~�9t 2145t 75pw        sq ~�ί�z[q ~ q ~�9t 2145t 84pw@@�鹙�sq ~�ί�v=q ~ q ~�9t 2146t 61pw        sq ~�ί�~q ~ q ~�9t 2146t 84pw@5oz�G�sq ~�ί�y�q ~ q ~�9t 2147t 61pw        sq ~�ίˁ�q ~ q ~�9t 2147t 84pw@5oz�G�sq ~�ίˁ�q ~ q ~�9t 2148t 75pw        sq ~�ί˅�q ~ q ~�9t 2148t 84pw@%�ʈ�sq ~�ίˁ�q ~ q ~�9t 2149t 61pw        sq ~�ίˉ_q ~ q ~�9t 2149t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 215t 75pw        sq ~��Z��q ~ q ~�9t 215t 84pw@5oz�G�sq ~�ί��Sq ~ q ~�9t 2150t 75pw        sq ~�ί���q ~ q ~�9t 2150t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2151t 61pw        sq ~�ί�߶q ~ q ~�9t 2151t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2152t 75pw        sq ~�ί��wq ~ q ~�9t 2152t 84pw@M]��%��sq ~�ί��Yq ~ q ~�9t 2153t 61pw        sq ~�ί��8q ~ q ~�9t 2153t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2154t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2155t 75pw        sq ~�ί��q ~ q ~�9t 2155t 84pw@$      sq ~�ί��q ~ q ~�9t 2156t 61pw        sq ~�ί��{q ~ q ~�9t 2156t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2157t 75pw        sq ~�ί��<q ~ q ~�9t 2157t 84pw@F�U�i�sq ~�ί��[q ~ q ~�9t 2158t 75pw        sq ~�ί���q ~ q ~�9t 2158t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2159t 61pw        sq ~�ί���q ~ q ~�9t 2159t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 216t 61pw        sq ~��Z��rq ~ q ~�9t 216t 84pw@5oz�G�sq ~�ί�L�q ~ q ~�9t 2160t 75pw        sq ~�ί�PTq ~ q ~�9t 2160t 84pw@@�鹙�sq ~�ί�Tq ~ q ~�9t 2161t 84pw@5oz�G�sq ~�ί�T4q ~ q ~�9t 2162t 75pw        sq ~�ί�W�q ~ q ~�9t 2162t 84pw@5oz�G�sq ~�ί�W�q ~ q ~�9t 2163t 75pw        sq ~�ί�[�q ~ q ~�9t 2163t 84pw@$      sq ~�ί�_Xq ~ q ~�9t 2164t 84pw@5oz�G�sq ~�ί�cq ~ q ~�9t 2165t 84pw@5oz�G�sq ~�ί�c8q ~ q ~�9t 2166t 75pw        sq ~�ί�f�q ~ q ~�9t 2166t 84pw@@�鹙�sq ~�ί�b�q ~ q ~�9t 2167t 61pw        sq ~�ί�j�q ~ q ~�9t 2167t 84pw@$      sq ~�ί�j�q ~ q ~�9t 2168t 75pw        sq ~�ί�n\q ~ q ~�9t 2168t 84pw@5oz�G�sq ~�ί�rq ~ q ~�9t 2169t 84pw@5oz�G�sq ~��Z��Tq ~ q ~�9t 217t 61pw        sq ~��Z��3q ~ q ~�9t 217t 84pw@5oz�G�sq ~�ί�ĳq ~ q ~�9t 2170t 84pw@@�鹙�sq ~�ί��tq ~ q ~�9t 2171t 84pw@F�U�i�sq ~�ί��5q ~ q ~�9t 2172t 84pw@@�鹙�sq ~�ί��Tq ~ q ~�9t 2173t 75pw        sq ~�ί���q ~ q ~�9t 2173t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2174t 75pw        sq ~�ί�ӷq ~ q ~�9t 2174t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2175t 75pw        sq ~�ί��xq ~ q ~�9t 2175t 84pw@5oz�G�sq ~�ί�חq ~ q ~�9t 2176t 75pw        sq ~�ί��9q ~ q ~�9t 2176t 84pw@@�鹙�sq ~�ί��Xq ~ q ~�9t 2177t 75pw        sq ~�ί���q ~ q ~�9t 2177t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2178t 61pw        sq ~�ί��q ~ q ~�9t 2178t 84pw@5oz�G�sq ~�ί��|q ~ q ~�9t 2179t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 218t 84pw@5oz�G�sq ~�ί�13q ~ q ~�9t 2180t 61pw        sq ~�ί�9q ~ q ~�9t 2180t 84pw@F�U�i�sq ~�ί�91q ~ q ~�9t 2181t 75pw        sq ~�ί�<�q ~ q ~�9t 2181t 84pw@@�鹙�sq ~�ί�@�q ~ q ~�9t 2182t 84pw@F�U�i�sq ~�ί�@�q ~ q ~�9t 2183t 75pw        sq ~�ί�DUq ~ q ~�9t 2183t 84pw@5oz�G�sq ~�ί�Dtq ~ q ~�9t 2184t 75pw        sq ~�ί�Hq ~ q ~�9t 2184t 84pw@F�U�i�sq ~�ί�C�q ~ q ~�9t 2185t 61pw        sq ~�ί�K�q ~ q ~�9t 2185t 84pw@5oz�G�sq ~�ί�K�q ~ q ~�9t 2186t 75pw        sq ~�ί�O�q ~ q ~�9t 2186t 84pw@$      sq ~�ί�O�q ~ q ~�9t 2187t 75pw        sq ~�ί�SYq ~ q ~�9t 2187t 84pw@F�U�i�sq ~�ί�Sxq ~ q ~�9t 2188t 75pw        sq ~�ί�Wq ~ q ~�9t 2188t 84pw@5oz�G�sq ~�ί�R�q ~ q ~�9t 2189t 61pw        sq ~�ί�Z�q ~ q ~�9t 2189t 84pw@$      sq ~��Z��q ~ q ~�9t 219t 75pw        sq ~��Z���q ~ q ~�9t 219t 84pw@@�鹙�sq ~�ίͩ�q ~ q ~�9t 2190t 75pw        sq ~�ίͭqq ~ q ~�9t 2190t 84pw@5oz�G�sq ~�ίͱ2q ~ q ~�9t 2191t 84pw@5oz�G�sq ~�ίͱQq ~ q ~�9t 2192t 75pw        sq ~�ίʹ�q ~ q ~�9t 2192t 84pw@5oz�G�sq ~�ί͵q ~ q ~�9t 2193t 75pw        sq ~�ί͸�q ~ q ~�9t 2193t 84pw@$      sq ~�ίͼuq ~ q ~�9t 2194t 84pw@$      sq ~�ίͼ�q ~ q ~�9t 2195t 75pw        sq ~�ί��6q ~ q ~�9t 2195t 84pw@$      sq ~�ί���q ~ q ~�9t 2196t 84pw@5oz�G�sq ~�ί�Ǹq ~ q ~�9t 2197t 84pw@M]��%��sq ~�ί�Úq ~ q ~�9t 2198t 61pw        sq ~�ί��yq ~ q ~�9t 2198t 84pw@8��A�sq ~�ί�˘q ~ q ~�9t 2199t 75pw        sq ~�ί��:q ~ q ~�9t 2199t 84pw@5oz�G�sq ~��W���q ~ q ~�9t 22t 0pw�ً���sq ~��Wŝq ~ q ~�9t 22t 12pw��H�Y�	sq ~��Wŝ�q ~ q ~�9t 22t 18pw@4�j��� sq ~��WŤ�q ~ q ~�9t 22t 32pw��� ��sq ~��Wť3q ~ q ~�9t 22t 37pw��b�8)_�sq ~��WŨ�q ~ q ~�9t 22t 46pw��=��ósq ~��W��q ~ q ~�9t 22t 5pw        sq ~��Z�?lq ~ q ~�9t 220t 61pw        sq ~��Z�GKq ~ q ~�9t 220t 84pw@5oz�G�sq ~�ίץ�q ~ q ~�9t 2200t 61pw        sq ~�ί׭�q ~ q ~�9t 2200t 84pw@5oz�G�sq ~�ί׭�q ~ q ~�9t 2201t 75pw        sq ~�ίױ\q ~ q ~�9t 2201t 84pw@5oz�G�sq ~�ί׭>q ~ q ~�9t 2202t 61pw        sq ~�ί׵q ~ q ~�9t 2202t 84pw@5oz�G�sq ~�ί׸�q ~ q ~�9t 2203t 84pw@$      sq ~�ί׼�q ~ q ~�9t 2204t 84pw@@�鹙�sq ~�ί׸�q ~ q ~�9t 2205t 61pw        sq ~�ί��`q ~ q ~�9t 2205t 84pw@5oz�G�sq ~�ί��!q ~ q ~�9t 2206t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2207t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2208t 61pw�������sq ~�ί�ˣq ~ q ~�9t 2208t 84pw@%��rBsq ~�ί�ǅq ~ q ~�9t 2209t 61pw        sq ~�ί��dq ~ q ~�9t 2209t 84pw@5oz�G�sq ~��Z�C-q ~ q ~�9t 221t 61pw        sq ~��Z�Kq ~ q ~�9t 221t 84pw@5oz�G�sq ~�ί�Xq ~ q ~�9t 2210t 75pw        sq ~�ί�!�q ~ q ~�9t 2210t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2211t 61pw        sq ~�ί�%�q ~ q ~�9t 2211t 84pw@@�鹙�sq ~�ί�%�q ~ q ~�9t 2212t 75pw        sq ~�ί�)|q ~ q ~�9t 2212t 84pw@#�hr�Nsq ~�ί�-=q ~ q ~�9t 2213t 84pw@5oz�G�sq ~�ί�)q ~ q ~�9t 2214t 61pw        sq ~�ί�0�q ~ q ~�9t 2214t 84pw@$      sq ~�ί�,�q ~ q ~�9t 2215t 61pw        sq ~�ί�4�q ~ q ~�9t 2215t 84pw@@�鹙�sq ~�ί�4�q ~ q ~�9t 2216t 75pw        sq ~�ί�8�q ~ q ~�9t 2216t 84pw@5oz�G�sq ~�ί�8�q ~ q ~�9t 2217t 75pw        sq ~�ί�<Aq ~ q ~�9t 2217t 84pw@5oz�G�sq ~�ί�8#q ~ q ~�9t 2218t 61pw        sq ~�ί�@q ~ q ~�9t 2218t 84pw@5oz�G�sq ~�ί�@!q ~ q ~�9t 2219t 75pw        sq ~�ί�C�q ~ q ~�9t 2219t 84pw@@�鹙�sq ~��Z�F�q ~ q ~�9t 222t 61pw        sq ~��Z�N�q ~ q ~�9t 222t 84pw@$      sq ~�ίؒ�q ~ q ~�9t 2220t 75pw        sq ~�ίؖYq ~ q ~�9t 2220t 84pw@5oz�G�sq ~�ίؖxq ~ q ~�9t 2221t 75pw        sq ~�ίؚq ~ q ~�9t 2221t 84pw@5oz�G�sq ~�ίؕ�q ~ q ~�9t 2222t 61pw        sq ~�ί؝�q ~ q ~�9t 2222t 84pw@5oz�G�sq ~�ίء�q ~ q ~�9t 2223t 84pw@5oz�G�sq ~�ίإ]q ~ q ~�9t 2224t 84pw@5oz�G�sq ~�ίةq ~ q ~�9t 2225t 84pw@$      sq ~�ίج�q ~ q ~�9t 2226t 84pw@@�鹙�sq ~�ίج�q ~ q ~�9t 2227t 75pw        sq ~�ίذ�q ~ q ~�9t 2227t 84pw@$      sq ~�ίشaq ~ q ~�9t 2228t 84pw@@�鹙�sq ~�ίش�q ~ q ~�9t 2229t 75pw        sq ~�ίظ"q ~ q ~�9t 2229t 84pw@5oz�G�sq ~��Z�N�q ~ q ~�9t 223t 75pw        sq ~��Z�R�q ~ q ~�9t 223t 84pw@$      sq ~�ί�
�q ~ q ~�9t 2230t 84pw@$      sq ~�ί�
�q ~ q ~�9t 2231t 75pw        sq ~�ί�yq ~ q ~�9t 2231t 84pw@@�鹙�sq ~�ί�
[q ~ q ~�9t 2232t 61pw        sq ~�ί�:q ~ q ~�9t 2232t 84pw@$      sq ~�ί�Yq ~ q ~�9t 2233t 75pw        sq ~�ί��q ~ q ~�9t 2233t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2234t 61pw        sq ~�ί��q ~ q ~�9t 2234t 84pw@$      sq ~�ί�}q ~ q ~�9t 2235t 84pw@@�鹙�sq ~�ί�!>q ~ q ~�9t 2236t 84pw@$      sq ~�ί�!]q ~ q ~�9t 2237t 75pw        sq ~�ί�$�q ~ q ~�9t 2237t 84pw@@�鹙�sq ~�ί� �q ~ q ~�9t 2238t 61pw        sq ~�ί�(�q ~ q ~�9t 2238t 84pw@F�U�i�sq ~�ί�,�q ~ q ~�9t 2239t 84pw@5oz�G�sq ~��Z�VOq ~ q ~�9t 224t 84pw@5oz�G�sq ~�ί�{uq ~ q ~�9t 2240t 75pw        sq ~�ί�q ~ q ~�9t 2240t 84pw@@�鹙�sq ~�ίق�q ~ q ~�9t 2241t 84pw@F�U�i�sq ~�ίق�q ~ q ~�9t 2242t 75pw        sq ~�ίن�q ~ q ~�9t 2242t 84pw@5oz�G�sq ~�ίيZq ~ q ~�9t 2243t 84pw@5oz�G�sq ~�ίَq ~ q ~�9t 2244t 84pw@5oz�G�sq ~�ίى�q ~ q ~�9t 2245t 61pw        sq ~�ίّ�q ~ q ~�9t 2245t 84pw@$      sq ~�ίٕ�q ~ q ~�9t 2246t 84pw@5oz�G�sq ~�ίٕ�q ~ q ~�9t 2247t 75pw        sq ~�ίٙ^q ~ q ~�9t 2247t 84pw@$      sq ~�ίٝq ~ q ~�9t 2248t 84pw@F�U�i�sq ~�ί٠�q ~ q ~�9t 2249t 84pw@5oz�G�sq ~��Z�R1q ~ q ~�9t 225t 61pw        sq ~��Z�Zq ~ q ~�9t 225t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2250t 61pw        sq ~�ί��vq ~ q ~�9t 2250t 84pw@5oz�G�sq ~�ί��7q ~ q ~�9t 2251t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2252t 61pw        sq ~�ί���q ~ q ~�9t 2252t 84pw@$      sq ~�ί���q ~ q ~�9t 2253t 84pw@5oz�G�sq ~�ί�zq ~ q ~�9t 2254t 84pw@5oz�G�sq ~�ί��\q ~ q ~�9t 2255t 61pw        sq ~�ί�;q ~ q ~�9t 2255t 84pw@$      sq ~�ί�	�q ~ q ~�9t 2256t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2257t 84pw@$      sq ~�ί��q ~ q ~�9t 2258t 75pw        sq ~�ί�~q ~ q ~�9t 2258t 84pw@@�鹙�sq ~�ί�?q ~ q ~�9t 2259t 84pw@5oz�G�sq ~��Z�U�q ~ q ~�9t 226t 61pw        sq ~��Z�]�q ~ q ~�9t 226t 84pw@5oz�G�sq ~�ί�d3q ~ q ~�9t 2260t 75pw        sq ~�ί�g�q ~ q ~�9t 2260t 84pw@@�鹙�sq ~�ί�c�q ~ q ~�9t 2261t 61pw        sq ~�ί�k�q ~ q ~�9t 2261t 84pw@5oz�G�sq ~�ί�k�q ~ q ~�9t 2262t 75pw        sq ~�ί�oWq ~ q ~�9t 2262t 84pw@'�����sq ~�ί�ovq ~ q ~�9t 2263t 75pw        sq ~�ί�sq ~ q ~�9t 2263t 84pw@5oz�G�sq ~�ί�v�q ~ q ~�9t 2264t 84pw@$      sq ~�ί�v�q ~ q ~�9t 2265t 75pw        sq ~�ί�z�q ~ q ~�9t 2265t 84pw@5oz�G�sq ~�ί�z�q ~ q ~�9t 2266t 75pw        sq ~�ί�~[q ~ q ~�9t 2266t 84pw@%��� ��sq ~�ίڂq ~ q ~�9t 2267t 84pw@5oz�G�sq ~�ίڂ;q ~ q ~�9t 2268t 75pw        sq ~�ίڅ�q ~ q ~�9t 2268t 84pw@@�鹙�sq ~�ίډ�q ~ q ~�9t 2269t 84pw@5oz�G�sq ~��Z�Y�q ~ q ~�9t 227t 61pw        sq ~��Z�a�q ~ q ~�9t 227t 84pw@@�鹙�sq ~�ί��4q ~ q ~�9t 2270t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2271t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2272t 61pw        sq ~�ί��q ~ q ~�9t 2272t 84pw@@�鹙�sq ~�ί�ߘq ~ q ~�9t 2273t 61pw        sq ~�ί��wq ~ q ~�9t 2273t 84pw@F�U�i�sq ~�ί��Yq ~ q ~�9t 2274t 61pw        sq ~�ί��8q ~ q ~�9t 2274t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2275t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2276t 61pw        sq ~�ί��q ~ q ~�9t 2276t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2277t 75pw        sq ~�ί��{q ~ q ~�9t 2277t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2278t 75pw        sq ~�ί��<q ~ q ~�9t 2278t 84pw@F�U�i�sq ~�ί��[q ~ q ~�9t 2279t 75pw        sq ~�ί���q ~ q ~�9t 2279t 84pw@$      sq ~��Z�]tq ~ q ~�9t 228t 61pw        sq ~��Z�eSq ~ q ~�9t 228t 84pw@@�鹙�sq ~�ί�P�q ~ q ~�9t 2280t 84pw@$      sq ~�ί�TTq ~ q ~�9t 2281t 84pw@5oz�G�sq ~�ί�Tsq ~ q ~�9t 2282t 75pw        sq ~�ί�Xq ~ q ~�9t 2282t 84pw@$      sq ~�ί�S�q ~ q ~�9t 2283t 61pw        sq ~�ί�[�q ~ q ~�9t 2283t 84pw@@�鹙�sq ~�ί�W�q ~ q ~�9t 2284t 61pw        sq ~�ί�_�q ~ q ~�9t 2284t 84pw@5oz�G�sq ~�ί�cXq ~ q ~�9t 2285t 84pw@5oz�G�sq ~�ί�cwq ~ q ~�9t 2286t 75pw        sq ~�ί�gq ~ q ~�9t 2286t 84pw@5oz�G�sq ~�ί�b�q ~ q ~�9t 2287t 61pw        sq ~�ί�j�q ~ q ~�9t 2287t 84pw@@�鹙�sq ~�ί�n�q ~ q ~�9t 2288t 84pw@$      sq ~�ί�j}q ~ q ~�9t 2289t 61pw        sq ~�ί�r\q ~ q ~�9t 2289t 84pw@@�鹙�sq ~��Z�a5q ~ q ~�9t 229t 61pw        sq ~��Z�iq ~ q ~�9t 229t 84pw@@�鹙�sq ~�ί��Pq ~ q ~�9t 2290t 75pw        sq ~�ί���q ~ q ~�9t 2290t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2291t 75pw        sq ~�ί�ȳq ~ q ~�9t 2291t 84pw@$      sq ~�ί��tq ~ q ~�9t 2292t 84pw@5oz�G�sq ~�ί��5q ~ q ~�9t 2293t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2294t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2295t 61pw        sq ~�ί�׷q ~ q ~�9t 2295t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2296t 75pw        sq ~�ί��xq ~ q ~�9t 2296t 84pw@5oz�G�sq ~�ί�ۗq ~ q ~�9t 2297t 75pw        sq ~�ί��9q ~ q ~�9t 2297t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2298t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2299t 75pw        sq ~�ί��q ~ q ~�9t 2299t 84pw@@�鹙�sq ~��WŠ�q ~ q ~�9t 23t 12pw?�5�K�0sq ~��WŤ�q ~ q ~�9t 23t 22pw����F�Osq ~��Wũq ~ q ~�9t 23t 38pw?��P�o�sq ~��Wũ2q ~ q ~�9t 23t 39pw@$      sq ~��Z���q ~ q ~�9t 230t 61pw        sq ~��Z���q ~ q ~�9t 230t 84pw@5oz�G�sq ~�ί��zq ~ q ~�9t 2300t 75pw        sq ~�ί��q ~ q ~�9t 2300t 84pw@5oz�G�sq ~�ί��;q ~ q ~�9t 2301t 75pw        sq ~�ί���q ~ q ~�9t 2301t 84pw@5oz�G�sq ~�ί�Ŀq ~ q ~�9t 2302t 61pw        sq ~�ί�̞q ~ q ~�9t 2302t 84pw@F�U�i�sq ~�ί�̽q ~ q ~�9t 2303t 75pw        sq ~�ί��_q ~ q ~�9t 2303t 84pw@5oz�G�sq ~�ί��~q ~ q ~�9t 2304t 75pw        sq ~�ί�� q ~ q ~�9t 2304t 84pw@$      sq ~�ί��q ~ q ~�9t 2305t 61pw        sq ~�ί���q ~ q ~�9t 2305t 84pw@$      sq ~�ί���q ~ q ~�9t 2306t 61pw        sq ~�ί�ۢq ~ q ~�9t 2306t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2307t 75pw        sq ~�ί��cq ~ q ~�9t 2307t 84pw@$      sq ~�ί��$q ~ q ~�9t 2308t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2309t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 231t 75pw        sq ~��Z��kq ~ q ~�9t 231t 84pw@F�U�i�sq ~�ί�1�q ~ q ~�9t 2310t 61pw        sq ~�ί�9{q ~ q ~�9t 2310t 84pw@5oz�G�sq ~�ί�=<q ~ q ~�9t 2311t 84pw@5oz�G�sq ~�ί�=[q ~ q ~�9t 2312t 75pw        sq ~�ί�@�q ~ q ~�9t 2312t 84pw@5oz�G�sq ~�ί�Aq ~ q ~�9t 2313t 75pw        sq ~�ί�D�q ~ q ~�9t 2313t 84pw@$      sq ~�ί�D�q ~ q ~�9t 2314t 75pw        sq ~�ί�Hq ~ q ~�9t 2314t 84pw@5oz�G�sq ~�ί�H�q ~ q ~�9t 2315t 75pw        sq ~�ί�L@q ~ q ~�9t 2315t 84pw@5oz�G�sq ~�ί�Pq ~ q ~�9t 2316t 84pw@@�鹙�sq ~�ί�K�q ~ q ~�9t 2317t 61pw        sq ~�ί�S�q ~ q ~�9t 2317t 84pw@$      sq ~�ί�S�q ~ q ~�9t 2318t 75pw        sq ~�ί�W�q ~ q ~�9t 2318t 84pw@$      sq ~�ί�[Dq ~ q ~�9t 2319t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 232t 75pw        sq ~��Z��,q ~ q ~�9t 232t 84pw@$      sq ~�ί��q ~ q ~�9t 2320t 61pw        sq ~�ί��q ~ q ~�9t 2320t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2321t 75pw        sq ~�ί汛q ~ q ~�9t 2321t 84pw@5oz�G�sq ~�ί�\q ~ q ~�9t 2322t 84pw@5oz�G�sq ~�ί�>q ~ q ~�9t 2323t 61pw        sq ~�ί�q ~ q ~�9t 2323t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2324t 61pw        sq ~�ί��q ~ q ~�9t 2324t 84pw@$      sq ~�ί��q ~ q ~�9t 2325t 61pw        sq ~�ί���q ~ q ~�9t 2325t 84pw@$      sq ~�ί���q ~ q ~�9t 2326t 75pw        sq ~�ί��`q ~ q ~�9t 2326t 84pw@5oz�G�sq ~�ί��!q ~ q ~�9t 2327t 84pw@@�鹙�sq ~�ί��@q ~ q ~�9t 2328t 75pw        sq ~�ί���q ~ q ~�9t 2328t 84pw@$7��O�sq ~�ί��q ~ q ~�9t 2329t 75pw        sq ~�ί�ϣq ~ q ~�9t 2329t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 233t 84pw@@�鹙�sq ~�ί�"9q ~ q ~�9t 2330t 84pw@@�鹙�sq ~�ί�%�q ~ q ~�9t 2331t 84pw@@�鹙�sq ~�ί�!�q ~ q ~�9t 2332t 61pw        sq ~�ί�)�q ~ q ~�9t 2332t 84pw@5oz�G�sq ~�ί�)�q ~ q ~�9t 2333t 75pw        sq ~�ί�-|q ~ q ~�9t 2333t 84pw@@�鹙�sq ~�ί�)^q ~ q ~�9t 2334t 61pw        sq ~�ί�1=q ~ q ~�9t 2334t 84pw@$      sq ~�ί�-q ~ q ~�9t 2335t 61pw        sq ~�ί�4�q ~ q ~�9t 2335t 84pw@$      sq ~�ί�5q ~ q ~�9t 2336t 75pw        sq ~�ί�8�q ~ q ~�9t 2336t 84pw@@�鹙�sq ~�ί�<�q ~ q ~�9t 2337t 84pw@@�鹙�sq ~�ί�<�q ~ q ~�9t 2338t 75pw        sq ~�ί�@Aq ~ q ~�9t 2338t 84pw@5oz�G�sq ~�ί�<#q ~ q ~�9t 2339t 61pw        sq ~�ί�Dq ~ q ~�9t 2339t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 234t 61pw        sq ~��Z�ʮq ~ q ~�9t 234t 84pw@@�鹙�sq ~�ί疘q ~ q ~�9t 2340t 84pw@@�鹙�sq ~�ί�zq ~ q ~�9t 2341t 61pw        sq ~�ί�Yq ~ q ~�9t 2341t 84pw@5oz�G�sq ~�ί�xq ~ q ~�9t 2342t 75pw        sq ~�ί�q ~ q ~�9t 2342t 84pw@$      sq ~�ί�9q ~ q ~�9t 2343t 75pw        sq ~�ί��q ~ q ~�9t 2343t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2344t 75pw        sq ~�ί祜q ~ q ~�9t 2344t 84pw@5oz�G�sq ~�ί�~q ~ q ~�9t 2345t 61pw        sq ~�ί�]q ~ q ~�9t 2345t 84pw@5oz�G�sq ~�ί�|q ~ q ~�9t 2346t 75pw        sq ~�ί�q ~ q ~�9t 2346t 84pw@M]��%��sq ~�ί� q ~ q ~�9t 2347t 61pw        sq ~�ί��q ~ q ~�9t 2347t 84pw@$      sq ~�ί素q ~ q ~�9t 2348t 84pw@@�鹙�sq ~�ί�aq ~ q ~�9t 2349t 84pw@5oz�G�sq ~��Z��oq ~ q ~�9t 235t 84pw@5oz�G�sq ~�ί�
�q ~ q ~�9t 2350t 84pw@$      sq ~�ί��q ~ q ~�9t 2351t 61pw        sq ~�ί��q ~ q ~�9t 2351t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2352t 75pw        sq ~�ί�yq ~ q ~�9t 2352t 84pw@5oz�G�sq ~�ί�:q ~ q ~�9t 2353t 84pw@5oz�G�sq ~�ί�Yq ~ q ~�9t 2354t 75pw        sq ~�ί��q ~ q ~�9t 2354t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2355t 61pw        sq ~�ί��q ~ q ~�9t 2355t 84pw@$      sq ~�ί��q ~ q ~�9t 2356t 61pw        sq ~�ί�!}q ~ q ~�9t 2356t 84pw@@�鹙�sq ~�ί�!�q ~ q ~�9t 2357t 75pw        sq ~�ί�%>q ~ q ~�9t 2357t 84pw@5oz�G�sq ~�ί�(�q ~ q ~�9t 2358t 84pw@5oz�G�sq ~�ί�,�q ~ q ~�9t 2359t 84pw@F�U�i�sq ~��Z�Ύq ~ q ~�9t 236t 75pw        sq ~��Z��0q ~ q ~�9t 236t 84pw@@�鹙�sq ~�ί�Vq ~ q ~�9t 2360t 84pw@5oz�G�sq ~�ί�q ~ q ~�9t 2361t 84pw@@�鹙�sq ~�ί�6q ~ q ~�9t 2362t 75pw        sq ~�ί��q ~ q ~�9t 2362t 84pw@$      sq ~�ί芙q ~ q ~�9t 2363t 84pw@5oz�G�sq ~�ί�Zq ~ q ~�9t 2364t 84pw@F�U�i�sq ~�ί�yq ~ q ~�9t 2365t 75pw        sq ~�ί�q ~ q ~�9t 2365t 84pw@F�U�i�sq ~�ί��q ~ q ~�9t 2366t 84pw@5oz�G�sq ~�ί虝q ~ q ~�9t 2367t 84pw@5oz�G�sq ~�ί�q ~ q ~�9t 2368t 61pw        sq ~�ί�^q ~ q ~�9t 2368t 84pw@5oz�G�sq ~�ί�@q ~ q ~�9t 2369t 61pw        sq ~�ί�q ~ q ~�9t 2369t 84pw@5oz�G�sq ~��Z��Oq ~ q ~�9t 237t 75pw        sq ~��Z���q ~ q ~�9t 237t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2370t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2371t 61pw        sq ~�ί��vq ~ q ~�9t 2371t 84pw@$      sq ~�ί��Xq ~ q ~�9t 2372t 61pw        sq ~�ί��7q ~ q ~�9t 2372t 84pw@@�鹙�sq ~�ί��Vq ~ q ~�9t 2373t 75pw        sq ~�ί���q ~ q ~�9t 2373t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2374t 61pw        sq ~�ί��q ~ q ~�9t 2374t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2375t 61pw        sq ~�ί�zq ~ q ~�9t 2375t 84pw@5oz�G�sq ~�ί�
;q ~ q ~�9t 2376t 84pw@$      sq ~�ί�
Zq ~ q ~�9t 2377t 75pw        sq ~�ί��q ~ q ~�9t 2377t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2378t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2379t 75pw        sq ~�ί�~q ~ q ~�9t 2379t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 238t 75pw        sq ~��Z�ٲq ~ q ~�9t 238t 84pw@5oz�G�sq ~�ί�drq ~ q ~�9t 2380t 75pw        sq ~�ί�hq ~ q ~�9t 2380t 84pw@@�鹙�sq ~�ί�h3q ~ q ~�9t 2381t 75pw        sq ~�ί�k�q ~ q ~�9t 2381t 84pw@#��o�"sq ~�ί�o�q ~ q ~�9t 2382t 84pw@F�U�i�sq ~�ί�kxq ~ q ~�9t 2383t 61pw        sq ~�ί�sWq ~ q ~�9t 2383t 84pw@$      sq ~�ί�svq ~ q ~�9t 2384t 75pw        sq ~�ί�wq ~ q ~�9t 2384t 84pw@@�鹙�sq ~�ί�z�q ~ q ~�9t 2385t 84pw@5oz�G�sq ~�ί�z�q ~ q ~�9t 2386t 75pw        sq ~�ί�~�q ~ q ~�9t 2386t 84pw@F�U�i�sq ~�ί�z|q ~ q ~�9t 2387t 61pw        sq ~�ί�[q ~ q ~�9t 2387t 84pw@$      sq ~�ί�zq ~ q ~�9t 2388t 75pw        sq ~�ί�q ~ q ~�9t 2388t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2389t 84pw@@�鹙�sq ~��Z�Քq ~ q ~�9t 239t 61pw        sq ~��Z��sq ~ q ~�9t 239t 84pw@$      sq ~�ί�Ԕq ~ q ~�9t 2390t 61pw        sq ~�ί��sq ~ q ~�9t 2390t 84pw@5oz�G�sq ~�ί�ܒq ~ q ~�9t 2391t 75pw        sq ~�ί��4q ~ q ~�9t 2391t 84pw@$      sq ~�ί���q ~ q ~�9t 2392t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2393t 75pw        sq ~�ί��q ~ q ~�9t 2393t 84pw@F�U�i�sq ~�ί��q ~ q ~�9t 2394t 61pw        sq ~�ί��wq ~ q ~�9t 2394t 84pw@$      sq ~�ί��Yq ~ q ~�9t 2395t 61pw        sq ~�ί��8q ~ q ~�9t 2395t 84pw@5oz�G�sq ~�ί��Wq ~ q ~�9t 2396t 75pw        sq ~�ί���q ~ q ~�9t 2396t 84pw@%�/�ͭ>sq ~�ί��q ~ q ~�9t 2397t 75pw        sq ~�ί���q ~ q ~�9t 2397t 84pw@$      sq ~�ί��{q ~ q ~�9t 2398t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2399t 75pw        sq ~�ί��<q ~ q ~�9t 2399t 84pw@@�鹙�sq ~��W��iq ~ q ~�9t 24t 0pw�"`��a+asq ~��WŤZq ~ q ~�9t 24t 10pw��)���>zsq ~��WŤ�q ~ q ~�9t 24t 12pw�
ƓJ��\sq ~��Wťq ~ q ~�9t 24t 16pw@%�p1Esq ~��WťRq ~ q ~�9t 24t 18pw@(����[�sq ~��WŨYq ~ q ~�9t 24t 22pw@�����sq ~��Wũq ~ q ~�9t 24t 28pw?ν�"sq ~��Wũ2q ~ q ~�9t 24t 29pw@)�~��C�sq ~��W���q ~ q ~�9t 24t 3pw��ϐ8Qsq ~��WŬ�q ~ q ~�9t 24t 37pw��X���K�sq ~��WŰWq ~ q ~�9t 24t 46pw@!��t�sq ~��W��q ~ q ~�9t 24t 5pw?�:���o�sq ~��Wų}q ~ q ~�9t 24t 51pw?�^"����sq ~��W��#q ~ q ~�9t 24t 6pw@'��)�Msq ~��W��Bq ~ q ~�9t 24t 7pw�����(�Gsq ~��Z�,gq ~ q ~�9t 240t 75pw        sq ~��Z�0	q ~ q ~�9t 240t 84pw@@�鹙�sq ~�ί�ܝq ~ q ~�9t 2400t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2401t 61pw        sq ~�ί��^q ~ q ~�9t 2401t 84pw@5oz�G�sq ~�ί��}q ~ q ~�9t 2402t 75pw        sq ~�ί��q ~ q ~�9t 2402t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2403t 84pw@$      sq ~�ί���q ~ q ~�9t 2404t 61pw        sq ~�ί��q ~ q ~�9t 2404t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2405t 61pw        sq ~�ί��bq ~ q ~�9t 2405t 84pw@@�鹙�sq ~�ί��Dq ~ q ~�9t 2406t 61pw        sq ~�ί��#q ~ q ~�9t 2406t 84pw@)�J
�sq ~�ί��Bq ~ q ~�9t 2407t 75pw        sq ~�ί���q ~ q ~�9t 2407t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2408t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2409t 61pw        sq ~�ί��fq ~ q ~�9t 2409t 84pw@$      sq ~��Z�3�q ~ q ~�9t 241t 84pw@$      sq ~�ί�MZq ~ q ~�9t 2410t 75pw        sq ~�ί�P�q ~ q ~�9t 2410t 84pw@@�鹙�sq ~�ί�L�q ~ q ~�9t 2411t 61pw        sq ~�ί�T�q ~ q ~�9t 2411t 84pw@@�鹙�sq ~�ί�P�q ~ q ~�9t 2412t 61pw        sq ~�ί�X~q ~ q ~�9t 2412t 84pw@5oz�G�sq ~�ί�X�q ~ q ~�9t 2413t 75pw        sq ~�ί�\?q ~ q ~�9t 2413t 84pw@'L�L��sq ~�ί�X!q ~ q ~�9t 2414t 61pw        sq ~�ί�` q ~ q ~�9t 2414t 84pw@@�鹙�sq ~�ί�[�q ~ q ~�9t 2415t 61pw        sq ~�ί�c�q ~ q ~�9t 2415t 84pw@5oz�G�sq ~�ί�_�q ~ q ~�9t 2416t 61pw        sq ~�ί�g�q ~ q ~�9t 2416t 84pw@5oz�G�sq ~�ί�g�q ~ q ~�9t 2417t 75pw        sq ~�ί�kCq ~ q ~�9t 2417t 84pw@$      sq ~�ί�kbq ~ q ~�9t 2418t 75pw        sq ~�ί�oq ~ q ~�9t 2418t 84pw@$      sq ~�ί�j�q ~ q ~�9t 2419t 61pw        sq ~�ί�r�q ~ q ~�9t 2419t 84pw@5oz�G�sq ~��Z�7�q ~ q ~�9t 242t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2420t 75pw        sq ~�ί��[q ~ q ~�9t 2420t 84pw@5oz�G�sq ~�ί��=q ~ q ~�9t 2421t 61pw        sq ~�ί��q ~ q ~�9t 2421t 84pw@$      sq ~�ί���q ~ q ~�9t 2422t 61pw        sq ~�ί���q ~ q ~�9t 2422t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2423t 75pw        sq ~�ί�Оq ~ q ~�9t 2423t 84pw@@�鹙�sq ~�ί�нq ~ q ~�9t 2424t 75pw        sq ~�ί��_q ~ q ~�9t 2424t 84pw@$      sq ~�ί��~q ~ q ~�9t 2425t 75pw        sq ~�ί�� q ~ q ~�9t 2425t 84pw@$      sq ~�ί��?q ~ q ~�9t 2426t 75pw        sq ~�ί���q ~ q ~�9t 2426t 84pw@$      sq ~�ί�� q ~ q ~�9t 2427t 75pw        sq ~�ί�ߢq ~ q ~�9t 2427t 84pw@@�鹙�sq ~�ί��cq ~ q ~�9t 2428t 84pw@5oz�G�sq ~�ί��$q ~ q ~�9t 2429t 84pw@%��Kߢ�sq ~��Z�7�q ~ q ~�9t 243t 75pw        sq ~��Z�;Lq ~ q ~�9t 243t 84pw@$      sq ~�ί�1�q ~ q ~�9t 2430t 61pw        sq ~�ί�9�q ~ q ~�9t 2430t 84pw@@�鹙�sq ~�ί�5�q ~ q ~�9t 2431t 61pw        sq ~�ί�={q ~ q ~�9t 2431t 84pw@5oz�G�sq ~�ί�=�q ~ q ~�9t 2432t 75pw        sq ~�ί�A<q ~ q ~�9t 2432t 84pw@5oz�G�sq ~�ί�=q ~ q ~�9t 2433t 61pw        sq ~�ί�D�q ~ q ~�9t 2433t 84pw@5oz�G�sq ~�ί�@�q ~ q ~�9t 2434t 61pw        sq ~�ί�H�q ~ q ~�9t 2434t 84pw@5oz�G�sq ~�ί�D�q ~ q ~�9t 2435t 61pw        sq ~�ί�Lq ~ q ~�9t 2435t 84pw@5oz�G�sq ~�ί�Haq ~ q ~�9t 2436t 61pw        sq ~�ί�P@q ~ q ~�9t 2436t 84pw@@�鹙�sq ~�ί�P_q ~ q ~�9t 2437t 75pw        sq ~�ί�Tq ~ q ~�9t 2437t 84pw@5oz�G�sq ~�ί�W�q ~ q ~�9t 2438t 84pw@@�鹙�sq ~�ί�W�q ~ q ~�9t 2439t 75pw        sq ~�ί�[�q ~ q ~�9t 2439t 84pw@5oz�G�sq ~��Z�?q ~ q ~�9t 244t 84pw@$      sq ~�ί��wq ~ q ~�9t 2440t 75pw        sq ~�ί��q ~ q ~�9t 2440t 84pw@$      sq ~�ί���q ~ q ~�9t 2441t 84pw@$      sq ~�ί���q ~ q ~�9t 2442t 75pw        sq ~�ί���q ~ q ~�9t 2442t 84pw@M]��%��sq ~�ί���q ~ q ~�9t 2443t 75pw        sq ~�ί��\q ~ q ~�9t 2443t 84pw@@�鹙�sq ~�ί��>q ~ q ~�9t 2444t 61pw        sq ~�ί��q ~ q ~�9t 2444t 84pw@@�鹙�sq ~�ί��<q ~ q ~�9t 2445t 75pw        sq ~�ί���q ~ q ~�9t 2445t 84pw@@�鹙�sq ~�ί�ğq ~ q ~�9t 2446t 84pw@5oz�G�sq ~�ί�ľq ~ q ~�9t 2447t 75pw        sq ~�ί��`q ~ q ~�9t 2447t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2448t 75pw        sq ~�ί��!q ~ q ~�9t 2448t 84pw@5oz�G�sq ~�ί��q ~ q ~�9t 2449t 61pw        sq ~�ί���q ~ q ~�9t 2449t 84pw@5oz�G�sq ~��Z�B�q ~ q ~�9t 245t 84pw@5oz�G�sq ~�ί�"xq ~ q ~�9t 2450t 84pw@5oz�G�sq ~�ί�&9q ~ q ~�9t 2451t 84pw@@�鹙�sq ~�ί�&Xq ~ q ~�9t 2452t 75pw        sq ~�ί�)�q ~ q ~�9t 2452t 84pw@@�鹙�sq ~�ί�%�q ~ q ~�9t 2453t 61pw        sq ~�ί�-�q ~ q ~�9t 2453t 84pw@F�U�i�sq ~�ί�)�q ~ q ~�9t 2454t 61pw        sq ~�ί�1|q ~ q ~�9t 2454t 84pw@F�U�i�sq ~�ί�1�q ~ q ~�9t 2455t 75pw        sq ~�ί�5=q ~ q ~�9t 2455t 84pw@5oz�G�sq ~�ί�8�q ~ q ~�9t 2456t 84pw@$      sq ~�ί�<�q ~ q ~�9t 2457t 84pw@@�鹙�sq ~�ί�<�q ~ q ~�9t 2458t 75pw        sq ~�ί�@�q ~ q ~�9t 2458t 84pw@5oz�G�sq ~�ί�@�q ~ q ~�9t 2459t 75pw        sq ~�ί�DAq ~ q ~�9t 2459t 84pw@&��]8�sq ~��Z�B�q ~ q ~�9t 246t 75pw        sq ~��Z�F�q ~ q ~�9t 246t 84pw@5oz�G�sq ~�ί��5q ~ q ~�9t 2460t 75pw        sq ~�ί���q ~ q ~�9t 2460t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2461t 61pw        sq ~�ί���q ~ q ~�9t 2461t 84pw@5oz�G�sq ~�ί��Yq ~ q ~�9t 2462t 84pw@$      sq ~�ί��q ~ q ~�9t 2463t 84pw@$      sq ~�ί���q ~ q ~�9t 2464t 84pw@5oz�G�sq ~�ί���q ~ q ~�9t 2465t 75pw        sq ~�ί���q ~ q ~�9t 2465t 84pw@$      sq ~�ί���q ~ q ~�9t 2466t 75pw        sq ~�ί��]q ~ q ~�9t 2466t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2467t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2468t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2469t 61pw        sq ~�ί���q ~ q ~�9t 2469t 84pw@$      sq ~��Z�Bqq ~ q ~�9t 247t 61pw        sq ~��Z�JPq ~ q ~�9t 247t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2470t 75pw        sq ~�ί�6q ~ q ~�9t 2470t 84pw@5oz�G�sq ~�ί�Uq ~ q ~�9t 2471t 75pw        sq ~�ί��q ~ q ~�9t 2471t 84pw@%����\sq ~�ί�
�q ~ q ~�9t 2472t 61pw        sq ~�ί��q ~ q ~�9t 2472t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2473t 75pw        sq ~�ί�yq ~ q ~�9t 2473t 84pw@$      sq ~�ί�[q ~ q ~�9t 2474t 61pw        sq ~�ί�:q ~ q ~�9t 2474t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2475t 84pw@5oz�G�sq ~�ί�q ~ q ~�9t 2476t 75pw        sq ~�ί�!�q ~ q ~�9t 2476t 84pw@@�鹙�sq ~�ί�%}q ~ q ~�9t 2477t 84pw@5oz�G�sq ~�ί�)>q ~ q ~�9t 2478t 84pw@F�U�i�sq ~�ί�,�q ~ q ~�9t 2479t 84pw@@�鹙�sq ~��Z�F2q ~ q ~�9t 248t 61pw        sq ~��Z�Nq ~ q ~�9t 248t 84pw@$      sq ~�ί��q ~ q ~�9t 2480t 84pw@@�鹙�sq ~�ί��Vq ~ q ~�9t 2481t 84pw@@�鹙�sq ~�ί��q ~ q ~�9t 2482t 84pw@@�鹙�sq ~�ί���q ~ q ~�9t 2483t 84pw@$      sq ~�ί���q ~ q ~�9t 2484t 84pw@F�U�i�sq ~�ί���q ~ q ~�9t 2485t 75pw        sq ~�ί��Zq ~ q ~�9t 2485t 84pw@F�U�i�sq ~�ί��gq ~ q ~�9t 2486t 0pw?���;�=sq ~�ί�{�q ~ q ~�9t 2486t 12pw���9�3sq ~�ί�|Pq ~ q ~�9t 2486t 18pw���B�Esq ~�ί��!q ~ q ~�9t 2486t 6pw@���^>�sq ~�ί���q ~ q ~�9t 2487t 27pw?���/�B�sq ~�ί���q ~ q ~�9t 2488t 16pw���ϔ=sq ~�ί���q ~ q ~�9t 2488t 28pw?������sq ~�ί��Fq ~ q ~�9t 2488t 3pw@��K�A;sq ~�ί���q ~ q ~�9t 2488t 32pw@�z�ѣ�sq ~�ί��sq ~ q ~�9t 2488t 39pw        sq ~�ί���q ~ q ~�9t 2488t 46pw����J<�sq ~�ί��{q ~ q ~�9t 2489t 21pw?������sq ~�ί���q ~ q ~�9t 2489t 59pw        sq ~��Z�I�q ~ q ~�9t 249t 61pw        sq ~��Z�Q�q ~ q ~�9t 249t 84pw@F�U�i�sq ~�ί��nq ~ q ~�9t 2490t 24pw���<�Tsq ~�ί���q ~ q ~�9t 2490t 31pw@t4�I$Nsq ~�ί��sq ~ q ~�9t 2490t 52pw        sq ~�ί���q ~ q ~�9t 2490t 67pw��$�rz�sq ~�ί�% q ~ q ~�9t 2491t 1pw@�X�S3sq ~�ί�(�q ~ q ~�9t 2492t 0pw�jN�����sq ~�ί��q ~ q ~�9t 2492t 22pw?�
Iý8sq ~�ί��q ~ q ~�9t 2492t 37pw        sq ~�ί��q ~ q ~�9t 2493t 27pw@��ٷ�sq ~�ί��1q ~ q ~�9t 2493t 68pw���U��/Xsq ~�ί�0Dq ~ q ~�9t 2494t 0pw�~�6��zsq ~�ί��4q ~ q ~�9t 2494t 22pw?�gG��sq ~�ί��q ~ q ~�9t 2494t 38pw        sq ~�ί��q ~ q ~�9t 2495t 27pw@!�$�!|sq ~�ί��Qq ~ q ~�9t 2496t 27pw@���?�sq ~�ί�|q ~ q ~�9t 2496t 60pw        sq ~�ί���q ~ q ~�9t 2497t 24pw?�n�śv�sq ~�ί��q ~ q ~�9t 2497t 31pw���C���sq ~�ί�q ~ q ~�9t 2497t 67pw��E��"Ssq ~�ί�
q ~ q ~�9t 2497t 71pw        sq ~�ί�?Hq ~ q ~�9t 2498t 0pw�cE
���sq ~�ί��wq ~ q ~�9t 2498t 12pw@�͘,_sq ~�ί���q ~ q ~�9t 2498t 16pw�ݠ[D���sq ~�ί��1q ~ q ~�9t 2498t 18pw�T�l�?sq ~�ί���q ~ q ~�9t 2498t 32pw��P�a��sq ~�ί�6q ~ q ~�9t 2498t 46pw��S NPl�sq ~�ί�@!q ~ q ~�9t 2498t 7pw        sq ~�ί�C	q ~ q ~�9t 2499t 0pw@`���usq ~�ί��8q ~ q ~�9t 2499t 12pw@� F�ΰsq ~�ί���q ~ q ~�9t 2499t 22pw��O�J��sq ~�ί�Cfq ~ q ~�9t 2499t 3pw��C�S� Ksq ~�ί��q ~ q ~�9t 2499t 32pw��*ʐ� Esq ~�ί�tq ~ q ~�9t 2499t 38pw@"΃;��sq ~�ί��q ~ q ~�9t 2499t 39pw?�/,0�sq ~�ί��q ~ q ~�9t 2499t 46pw�����iGsq ~�ί�C�q ~ q ~�9t 2499t 5pw?��VQ�usq ~�ί�C�q ~ q ~�9t 2499t 6pw?��8e� �sq ~��WŨxq ~ q ~�9t 25t 13pw� �3Tsq ~��Wū�q ~ q ~�9t 25t 21pw@$      sq ~��WŬ�q ~ q ~�9t 25t 26pw@7��=��sq ~��W��q ~ q ~�9t 25t 4pw        sq ~��Wų�q ~ q ~�9t 25t 45pw� i�oe,�sq ~��Z���q ~ q ~�9t 250t 61pw        sq ~��Z��hq ~ q ~�9t 250t 84pw@@�鹙�sq ~�ΰ!jq ~ q ~�9t 2500t 0pw�H\ۅ�?sq ~�ΰٙq ~ q ~�9t 2500t 12pw@i;�Ǟsq ~�ΰ�q ~ q ~�9t 2500t 16pw�͏���5sq ~�ΰ�Zq ~ q ~�9t 2500t 22pw��jb��:*sq ~�ΰ�q ~ q ~�9t 2500t 28pw�ѳ�%��sq ~�ΰ�q ~ q ~�9t 2500t 32pw���M$�sq ~�ΰ��q ~ q ~�9t 2500t 39pw        sq ~�ΰ�Xq ~ q ~�9t 2500t 46pw����=sq ~�ΰ�Yq ~ q ~�9t 2501t 24pw?�L��Ҿ/sq ~�ΰ�9q ~ q ~�9t 2501t 35pw        sq ~�ΰ�q ~ q ~�9t 2502t 24pw@
ЬM�esq ~�ΰ�~q ~ q ~�9t 2502t 31pw��;�3z�sq ~�ΰ��q ~ q ~�9t 2502t 35pw���{~�u>sq ~�ΰ�q ~ q ~�9t 2502t 52pw���{~�u>sq ~�ΰ�>q ~ q ~�9t 2502t 53pw@�@��sq ~�ΰ�{q ~ q ~�9t 2502t 67pw��[��y�Csq ~�ΰ�8q ~ q ~�9t 2503t 27pw?��G��sq ~�ΰ�[q ~ q ~�9t 2503t 68pw        sq ~�ΰ��q ~ q ~�9t 2504t 49pw?�@�`e��sq ~�ΰ�#q ~ q ~�9t 2504t 72pw        sq ~�ΰ�=q ~ q ~�9t 2505t 35pw?�@�`e��sq ~�ΰ�bq ~ q ~�9t 2505t 52pw?�@�`e��sq ~�ΰ
(q ~ q ~�9t 2506t 80pw?�@�`e��sq ~�ΰ
�q ~ q ~�9t 2506t 83pw?�@�`e��sq ~�ΰ�q ~ q ~�9t 2507t 64pw?�@�`e��sq ~�ΰ�q ~ q ~�9t 2508t 48pw?�@�`e��sq ~�ΰ�bq ~ q ~�9t 2509t 12pw?�Xs��^sq ~�ΰ
(q ~ q ~�9t 2509t 50pw        sq ~��Z���q ~ q ~�9t 251t 75pw        sq ~��Z��)q ~ q ~�9t 251t 84pw@F�U�i�sq ~�ΰM�q ~ q ~�9t 2510t 12pw        sq ~�ΰ�&q ~ q ~�9t 2510t 3pw��=�Eܶsq ~�ΰV4q ~ q ~�9t 2510t 38pw?��f�sq ~�ΰY�q ~ q ~�9t 2510t 47pw@m�D�sq ~�ΰ��q ~ q ~�9t 2511t 0pw�	���sq ~�ΰQ�q ~ q ~�9t 2511t 12pw?�!=��!�sq ~�ΰUzq ~ q ~�9t 2511t 22pw@}�+��sq ~�ΰU�q ~ q ~�9t 2511t 23pw?u�ɏ;�sq ~�ΰV4q ~ q ~�9t 2511t 28pw?�[�|�a<sq ~�ΰVSq ~ q ~�9t 2511t 29pw?�s��Qr�sq ~�ΰ��q ~ q ~�9t 2511t 3pw��N�'�;sq ~�ΰY;q ~ q ~�9t 2511t 32pw@ ��RM-{sq ~�ΰY�q ~ q ~�9t 2511t 37pw        sq ~�ΰY�q ~ q ~�9t 2511t 38pw?�G�k<�sq ~�ΰ]�q ~ q ~�9t 2511t 47pw@J�lsq ~�ΰ�Kq ~ q ~�9t 2512t 0pw�����n�Gsq ~�ΰU<q ~ q ~�9t 2512t 10pw        sq ~�ΰY;q ~ q ~�9t 2512t 22pw��
�2f��sq ~�ΰaXq ~ q ~�9t 2512t 47pw@��(�%{sq ~�ΰYyq ~ q ~�9t 2513t 14pw@�O���sq ~�ΰY�q ~ q ~�9t 2513t 15pw���\pL�sq ~�ΰo�q ~ q ~�9t 2513t 72pw�3�_���sq ~�ΰ�q ~ q ~�9t 2513t 8pw@�h1z:sq ~�ΰ�#q ~ q ~�9t 2513t 9pw� >|>a7sq ~�ΰo�q ~ q ~�9t 2514t 61pw��K����Ysq ~�ΰw�q ~ q ~�9t 2514t 84pw@�n� =sq ~�ΰ`�q ~ q ~�9t 2515t 14pw@�%g�l�sq ~�ΰaq ~ q ~�9t 2515t 15pw��IЯw�;sq ~�ΰlq ~ q ~�9t 2515t 43pw        sq ~�ΰwCq ~ q ~�9t 2515t 72pw���H��Xsq ~�ΰ��q ~ q ~�9t 2515t 8pw�ˋA*#�sq ~�ΰ��q ~ q ~�9t 2515t 9pw�̮�]�sq ~�ΰ�Oq ~ q ~�9t 2516t 0pw�c��F� �sq ~�ΰe8q ~ q ~�9t 2516t 18pw�+Hf0ֹsq ~�ΰh�q ~ q ~�9t 2516t 28pw        sq ~�ΰ��q ~ q ~�9t 2516t 5pw?�\*��z-sq ~�ΰ�	q ~ q ~�9t 2516t 6pw@
-�_"8�sq ~�ΰ�q ~ q ~�9t 2517t 0pw��!	�\�sq ~�ΰh?q ~ q ~�9t 2517t 12pw?�Y���sq ~�ΰl q ~ q ~�9t 2517t 22pw@
$��w�Ysq ~�ΰ��q ~ q ~�9t 2517t 5pw?��E��CXsq ~�ΰ��q ~ q ~�9t 2517t 6pw?�0�6�gsq ~�ΰp\q ~ q ~�9t 2518t 27pw?��O�blsq ~�ΰs�q ~ q ~�9t 2519t 25pw@�GD��sq ~�ΰz�q ~ q ~�9t 2519t 40pw        sq ~��Z���q ~ q ~�9t 252t 84pw@5oz�G�sq ~�ΰ
(q ~ q ~�9t 2520t 0pw?�i��Rsq ~�ΰ�Wq ~ q ~�9t 2520t 12pw?�KAI1�sq ~�ΰ��q ~ q ~�9t 2520t 29pw        sq ~�ΰƔq ~ q ~�9t 2521t 16pw?��u9�	�sq ~�ΰ��q ~ q ~�9t 2521t 46pw?���s��sq ~�ΰ��q ~ q ~�9t 2521t 47pw�Xc� �xksq ~�ΰ��q ~ q ~�9t 2521t 50pw        sq ~�ΰ��q ~ q ~�9t 2522t 12pw��m8E��sq ~�ΰʓq ~ q ~�9t 2522t 18pw        sq ~�ΰ͚q ~ q ~�9t 2522t 22pw���j�9�sq ~�ΰ�Tq ~ q ~�9t 2522t 28pw���l����sq ~�ΰ�[q ~ q ~�9t 2522t 32pw����P�sq ~�ΰշq ~ q ~�9t 2522t 47pw�l^�-
<sq ~�ΰ�Tq ~ q ~�9t 2523t 18pw        sq ~�ΰ�q ~ q ~�9t 2523t 28pw?��j�sq ~�ΰ,q ~ q ~�9t 2524t 0pw        sq ~�ΰ��q ~ q ~�9t 2524t 32pw?Ķ�s
� sq ~�ΰ�q ~ q ~�9t 2524t 46pw?�C�9W.sq ~�ΰ�Zq ~ q ~�9t 2525t 14pw?��|�!�sq ~�ΰ�yq ~ q ~�9t 2525t 15pw��}A�p�	sq ~�ΰ�q ~ q ~�9t 2525t 72pw�dBrRF;ssq ~�ΰ�q ~ q ~�9t 2525t 8pw?žF[�Ssq ~�ΰq ~ q ~�9t 2525t 9pw�d���A_sq ~�ΰ�q ~ q ~�9t 2526t 14pw?��D����sq ~�ΰ�:q ~ q ~�9t 2526t 15pw��I���sq ~�ΰ�q ~ q ~�9t 2526t 41pw        sq ~�ΰ�cq ~ q ~�9t 2526t 72pw�և�Pb�sq ~�ΰ!�q ~ q ~�9t 2526t 8pw?�"ƴI�msq ~�ΰ!�q ~ q ~�9t 2526t 9pw��S!��/sq ~�ΰ��q ~ q ~�9t 2527t 14pw?�E����sq ~�ΰ��q ~ q ~�9t 2527t 15pw�ʩ�+!�;sq ~�ΰ� q ~ q ~�9t 2527t 43pw        sq ~�ΰ��q ~ q ~�9t 2528t 14pw@�_�Nsq ~�ΰ�q ~ q ~�9t 2528t 15pw�0*�oxsq ~�ΰ��q ~ q ~�9t 2528t 43pw        sq ~�ΰ��q ~ q ~�9t 2528t 72pw����f&�sq ~�ΰ)(q ~ q ~�9t 2528t 8pw?��`=�Bsq ~�ΰ)Gq ~ q ~�9t 2528t 9pw�����Vsq ~�ΰ�q ~ q ~�9t 2529t 24pw?�ݼ���Nsq ~�ΰ�Cq ~ q ~�9t 2529t 53pw        sq ~��Z��	q ~ q ~�9t 253t 75pw        sq ~��Z���q ~ q ~�9t 253t 84pw@$      sq ~�ΰ~�q ~ q ~�9t 2530t 0pw��^n�sq ~�ΰ:wq ~ q ~�9t 2530t 22pw?�K�i��lsq ~�ΰE|q ~ q ~�9t 2530t 50pw        sq ~�ΰ:�q ~ q ~�9t 2531t 14pw?����=sq ~�ΰ:�q ~ q ~�9t 2531t 15pw���N�P�sq ~�ΰ=�q ~ q ~�9t 2531t 20pw        sq ~�ΰP�q ~ q ~�9t 2531t 72pw���>�#�sq ~�ΰ�@q ~ q ~�9t 2531t 8pw?�J�'��Osq ~�ΰ�_q ~ q ~�9t 2531t 9pw��4 	N5�sq ~�ΰ�	q ~ q ~�9t 2532t 0pw���K��sq ~�ΰ>8q ~ q ~�9t 2532t 12pw?��N*�F~sq ~�ΰA�q ~ q ~�9t 2532t 22pw@���$�9sq ~�ΰB�q ~ q ~�9t 2532t 29pw        sq ~�ΰ��q ~ q ~�9t 2532t 6pw?��C�9�0sq ~�ΰB7q ~ q ~�9t 2533t 14pw@t!�D�sq ~�ΰBVq ~ q ~�9t 2533t 15pw��G��sq ~�ΰM[q ~ q ~�9t 2533t 43pw��8!Jsq ~�ΰNq ~ q ~�9t 2533t 49pw        sq ~�ΰXq ~ q ~�9t 2533t 72pw���V�OVsq ~�ΰ��q ~ q ~�9t 2533t 8pw?�3g���sq ~�ΰ��q ~ q ~�9t 2533t 9pw�����(0sq ~�ΰI�q ~ q ~�9t 2534t 24pw��*b��sq ~�ΰMq ~ q ~�9t 2534t 31pw��s�o�sq ~�ΰT�q ~ q ~�9t 2534t 54pw?���Q16Vsq ~�ΰYq ~ q ~�9t 2534t 67pw��!�̈sq ~�ΰMzq ~ q ~�9t 2535t 24pw@h��Hsq ~�ΰP�q ~ q ~�9t 2535t 31pw��݀�f�sq ~�ΰX�q ~ q ~�9t 2535t 54pw@\��r|sq ~�ΰ\�q ~ q ~�9t 2535t 67pw��q;a8�sq ~�ΰ_�q ~ q ~�9t 2535t 71pw        sq ~�ΰ_�q ~ q ~�9t 2536t 61pw        sq ~�ΰg�q ~ q ~�9t 2536t 84pw@Ʋ'�)�sq ~�ΰP�q ~ q ~�9t 2537t 10pw        sq ~�ΰP�q ~ q ~�9t 2537t 12pw?��0�~��sq ~�ΰT�q ~ q ~�9t 2538t 12pw?�[C_�j�sq ~�ΰYXq ~ q ~�9t 2538t 29pw        sq ~�ΰXq ~ q ~�9t 2539t 12pw?�[C_�j�sq ~�ΰ�
q ~ q ~�9t 2539t 6pw        sq ~��Z���q ~ q ~�9t 254t 61pw        sq ~��Z��lq ~ q ~�9t 254t 84pw@$      sq ~�ΰ�q ~ q ~�9t 2540t 12pw?��0�~��sq ~�ΰ��q ~ q ~�9t 2540t 18pw        sq ~�ΰ��q ~ q ~�9t 2541t 24pw@��=��Zsq ~�ΰ��q ~ q ~�9t 2542t 27pw�����<ksq ~�ΰ�q ~ q ~�9t 2542t 60pw@'cB���Bsq ~�ΰ�q ~ q ~�9t 2542t 68pw��]�Q��sq ~�ΰ��q ~ q ~�9t 2543t 14pw��b}�U@-sq ~�ΰ��q ~ q ~�9t 2543t 15pw@t�mWf�sq ~�ΰ�|q ~ q ~�9t 2543t 41pw���l��sq ~�ΰ��q ~ q ~�9t 2543t 43pw�����I�sq ~�ΰ��q ~ q ~�9t 2543t 72pw��;�sp�sq ~�ΰ�!q ~ q ~�9t 2543t 8pw���T���Qsq ~�ΰ�@q ~ q ~�9t 2543t 9pw?�!�|C� sq ~�ΰ�=q ~ q ~�9t 2544t 41pw@�@��sq ~�ΰ�{q ~ q ~�9t 2544t 43pw        sq ~�ΰq ~ q ~�9t 2544t 9pw@cC�`�@sq ~�ΰ�6q ~ q ~�9t 2545t 27pw?�e
�`��sq ~�ΰ�Yq ~ q ~�9t 2545t 68pw        sq ~�ΰŚq ~ q ~�9t 2546t 24pw?�����sq ~�ΰоq ~ q ~�9t 2546t 53pw        sq ~�ΰ�[q ~ q ~�9t 2547t 24pw?�<�Ǯ�ksq ~�ΰ�[q ~ q ~�9t 2548t 14pw?��0�O�sq ~�ΰ�9q ~ q ~�9t 2548t 49pw        sq ~�ΰߣq ~ q ~�9t 2548t 72pw���%lYJGsq ~�ΰ�q ~ q ~�9t 2548t 8pw?�w�`P�sq ~�ΰ�q ~ q ~�9t 2549t 0pw��C�S� Msq ~�ΰ̠q ~ q ~�9t 2549t 10pw        sq ~�ΰ�q ~ q ~�9t 2549t 38pw?���_�6sq ~��Z���q ~ q ~�9t 255t 75pw        sq ~��Z��-q ~ q ~�9t 255t 84pw@@�鹙�sq ~�ΰgEq ~ q ~�9t 2550t 0pw����D��sq ~�ΰtq ~ q ~�9t 2550t 12pw����dI/sq ~�ΰ .q ~ q ~�9t 2550t 18pw@���Mp"sq ~�ΰ#5q ~ q ~�9t 2550t 22pw��(P��sq ~�ΰ'�q ~ q ~�9t 2550t 37pw        sq ~�ΰ'�q ~ q ~�9t 2550t 38pw?���DZ�sq ~�ΰ'4q ~ q ~�9t 2551t 24pw?ﴄ2�ssq ~�ΰ*�q ~ q ~�9t 2551t 31pw���:�V�sq ~�ΰ2Xq ~ q ~�9t 2551t 53pw        sq ~�ΰ6�q ~ q ~�9t 2551t 67pw��&ssq ~�ΰ*�q ~ q ~�9t 2552t 24pw@ ��4sq ~�ΰ:Vq ~ q ~�9t 2552t 67pw        sq ~�ΰr�q ~ q ~�9t 2553t 0pw���~f.sq ~�ΰ*yq ~ q ~�9t 2553t 10pw        sq ~�ΰ*�q ~ q ~�9t 2553t 12pw@y{�24�sq ~�ΰ.xq ~ q ~�9t 2553t 22pw���a'�sq ~�ΰ2�q ~ q ~�9t 2553t 38pw@=NT�psq ~�ΰ6�q ~ q ~�9t 2553t 47pw���Z�ف^sq ~�ΰ.:q ~ q ~�9t 2554t 10pw        sq ~�ΰ.xq ~ q ~�9t 2554t 12pw?�A�&�sq ~�ΰ29q ~ q ~�9t 2555t 12pw@թHmp�sq ~�ΰ5�q ~ q ~�9t 2555t 22pw        sq ~�ΰzgq ~ q ~�9t 2555t 3pw��s���sq ~�ΰ5�q ~ q ~�9t 2556t 12pw?�A�$�sq ~�ΰ9�q ~ q ~�9t 2557t 12pw� �KNpsq ~�ΰA�q ~ q ~�9t 2557t 37pw        sq ~�ΰA{q ~ q ~�9t 2558t 24pw?ΡO�ybRsq ~�ΰL�q ~ q ~�9t 2558t 53pw        sq ~�ΰE<q ~ q ~�9t 2559t 24pw?�%ԩ��sq ~�ΰPAq ~ q ~�9t 2559t 52pw        sq ~��Z��q ~ q ~�9t 256t 61pw        sq ~��Z���q ~ q ~�9t 256t 84pw@$      sq ~�ΰ��q ~ q ~�9t 2560t 24pw?��2O�*psq ~�ΰ�:q ~ q ~�9t 2560t 71pw        sq ~�ΰ��q ~ q ~�9t 2561t 24pw?�%ԩ��sq ~�ΰ��q ~ q ~�9t 2561t 53pw        sq ~�ΰ��q ~ q ~�9t 2562t 60pw        sq ~�ΰ��q ~ q ~�9t 2562t 68pw?�cy�q9\sq ~�ΰ�q ~ q ~�9t 2563t 24pw?�eDa��sq ~�ΰ�yq ~ q ~�9t 2563t 31pw��ˣV+sq ~�ΰ�Xq ~ q ~�9t 2563t 54pw?��*�}sq ~�ΰ�vq ~ q ~�9t 2563t 67pw����Osq ~�ΰ��q ~ q ~�9t 2564t 12pw?�<f����sq ~�ΰ�qq ~ q ~�9t 2564t 29pw        sq ~�ΰ�q ~ q ~�9t 2564t 38pw���ɣsq ~�ΰ�q ~ q ~�9t 2565t 1pw?��U��6�sq ~�ΰ�]q ~ q ~�9t 2565t 62pw        sq ~�ΰ�Yq ~ q ~�9t 2566t 12pw��'.~!:�sq ~�ΰ�q ~ q ~�9t 2566t 22pw?��D���sq ~�ΰ��q ~ q ~�9t 2566t 28pw��x!w��Asq ~�ΰ��q ~ q ~�9t 2566t 32pw���I)�}-sq ~�ΰ��q ~ q ~�9t 2566t 38pw?߭_���sq ~�ΰ�7q ~ q ~�9t 2566t 47pw��;�L�Ժsq ~�ΰ�>q ~ q ~�9t 2566t 51pw        sq ~�ΰ�q ~ q ~�9t 2567t 24pw?9�sq ~�ΰ��q ~ q ~�9t 2567t 35pw        sq ~�ΰ�7q ~ q ~�9t 2568t 27pw?��=��sq ~�ΰ��q ~ q ~�9t 2569t 1pw?���v�sq ~�ΰ�aq ~ q ~�9t 2569t 62pw        sq ~��Z���q ~ q ~�9t 257t 61pw        sq ~��Z���q ~ q ~�9t 257t 84pw@@�鹙�sq ~�ΰ�q ~ q ~�9t 2570t 27pw?���v�sq ~�ΰ�q ~ q ~�9t 2571t 12pw?��"/^v�sq ~�ΰoq ~ q ~�9t 2571t 16pw����L�sq ~�ΰnq ~ q ~�9t 2571t 28pw��V�V� zsq ~�ΰT~q ~ q ~�9t 2571t 6pw        sq ~�ΰW�q ~ q ~�9t 2572t 0pw        sq ~�ΰ�q ~ q ~�9t 2572t 12pw@
` ��sq ~�ΰuq ~ q ~�9t 2573t 12pw?��"/^w�sq ~�ΰ�q ~ q ~�9t 2573t 28pw��˧�!�sq ~�ΰ\q ~ q ~�9t 2573t 7pw        sq ~�ΰ_&q ~ q ~�9t 2574t 1pw���I���sq ~�ΰ)�q ~ q ~�9t 2574t 62pw        sq ~�ΰSq ~ q ~�9t 2575t 27pw@#�r�͚sq ~�ΰ-~q ~ q ~�9t 2575t 60pw        sq ~�ΰ"�q ~ q ~�9t 2576t 24pw?��4-iqsq ~�ΰ&�q ~ q ~�9t 2576t 35pw��B5!@��sq ~�ΰ-�q ~ q ~�9t 2576t 52pw��B5!@��sq ~�ΰ-�q ~ q ~�9t 2576t 54pw@��߯�sq ~�ΰ"�q ~ q ~�9t 2577t 14pw?�n�qHsq ~�ΰ"�q ~ q ~�9t 2577t 15pw����P6�Gsq ~�ΰ-�q ~ q ~�9t 2577t 41pw        sq ~�ΰ-�q ~ q ~�9t 2578t 32pw?�m����sq ~�ΰ5 q ~ q ~�9t 2578t 50pw        sq ~�ΰ*9q ~ q ~�9t 2579t 14pw���+㕂nsq ~�ΰ*Xq ~ q ~�9t 2579t 15pw?��*/�sq ~�ΰ5]q ~ q ~�9t 2579t 43pw        sq ~�ΰ@�q ~ q ~�9t 2579t 72pw��9N�<sq ~�ΰr�q ~ q ~�9t 2579t 8pw��q Y?�ssq ~�ΰr�q ~ q ~�9t 2579t 9pw?��4v}�}sq ~��Z���q ~ q ~�9t 258t 75pw        sq ~��Z��pq ~ q ~�9t 258t 84pw@$      sq ~�ΰ|�q ~ q ~�9t 2580t 12pw?�h]sq ~�ΰ�qq ~ q ~�9t 2580t 23pw        sq ~�ΰ��q ~ q ~�9t 2581t 84pw?�h]sq ~�ΰ�q ~ q ~�9t 2582t 1pw@6���sq ~�ΰ�Tq ~ q ~�9t 2582t 66pw        sq ~�ΰ�0q ~ q ~�9t 2583t 27pw@oY,�sq ~�ΰ�Sq ~ q ~�9t 2583t 68pw        sq ~�ΰ�fq ~ q ~�9t 2584t 0pw���N�~Ksq ~�ΰ��q ~ q ~�9t 2584t 12pw?�]�ҕ�sq ~�ΰ�[q ~ q ~�9t 2584t 50pw        sq ~�ΰ��q ~ q ~�9t 2585t 61pw���N�8sq ~�ΰ��q ~ q ~�9t 2585t 84pw?�]�ҕ�sq ~�ΰ��q ~ q ~�9t 2586t 0pw�		q�H~sq ~�ΰ��q ~ q ~�9t 2586t 22pw@�ln��sq ~�ΰ�q ~ q ~�9t 2587t 14pw@����B�sq ~�ΰ�5q ~ q ~�9t 2587t 15pw���H����sq ~�ΰ�^q ~ q ~�9t 2587t 72pw��C����sq ~�ΰߡq ~ q ~�9t 2587t 8pw?���cR�	sq ~�ΰ��q ~ q ~�9t 2587t 9pw���zt\sq ~�ΰ��q ~ q ~�9t 2588t 24pw@I7͞��sq ~�ΰ��q ~ q ~�9t 2588t 31pw���	���sq ~�ΰ��q ~ q ~�9t 2588t 54pw        sq ~�ΰ��q ~ q ~�9t 2588t 67pw�����E�sq ~�ΰ�+q ~ q ~�9t 2589t 0pw�݀�2N�Rsq ~�ΰ�Zq ~ q ~�9t 2589t 12pw?�o�J�sq ~�ΰ��q ~ q ~�9t 2589t 6pw        sq ~��Z�q ~ q ~�9t 259t 75pw        sq ~��Z��1q ~ q ~�9t 259t 84pw@@�鹙�sq ~�ΰ�q ~ q ~�9t 2590t 61pw��D;�>sq ~�ΰ�q ~ q ~�9t 2590t 75pw        sq ~�ΰuq ~ q ~�9t 2590t 84pw?�o�J/sq ~�ΰ��q ~ q ~�9t 2591t 24pw?�N�Z�	sq ~�ΰ�q ~ q ~�9t 2591t 31pw��u�&)!sq ~�ΰ��q ~ q ~�9t 2591t 35pw���J(�T�sq ~�ΰ�q ~ q ~�9t 2591t 52pw���J(�T�sq ~�ΰ�q ~ q ~�9t 2591t 54pw        sq ~�ΰq ~ q ~�9t 2591t 67pw��2E!k&sq ~�ΰ@Cq ~ q ~�9t 2592t 0pw����#+:wsq ~�ΰ�4q ~ q ~�9t 2592t 10pw        sq ~�ΰ�rq ~ q ~�9t 2592t 12pw?�x֒6��sq ~�ΰ��q ~ q ~�9t 2592t 16pw��I��e�sq ~�ΰ�Rq ~ q ~�9t 2592t 23pw?���P��sq ~�ΰ��q ~ q ~�9t 2592t 28pw?���<��sq ~�ΰ�q ~ q ~�9t 2592t 29pw?���]l�sq ~�ΰ��q ~ q ~�9t 2592t 32pw?��{�}sq ~�ΰ �q ~ q ~�9t 2592t 37pw?�5�\��sq ~�ΰ1q ~ q ~�9t 2592t 46pw���v	��sq ~�ΰ�qq ~ q ~�9t 2593t 14pw@0�.��sq ~�ΰ��q ~ q ~�9t 2593t 15pw��� d��_sq ~�ΰOq ~ q ~�9t 2593t 49pw        sq ~�ΰ�q ~ q ~�9t 2593t 72pw��W����sq ~�ΰD�q ~ q ~�9t 2593t 8pw��oZf�&�sq ~�ΰEq ~ q ~�9t 2593t 9pw��!u�{1sq ~�ΰG�q ~ q ~�9t 2594t 0pw��ϐ8Tjsq ~�ΰ pq ~ q ~�9t 2594t 16pw?��}wC.sq ~�ΰ0q ~ q ~�9t 2594t 38pw        sq ~�ΰ�q ~ q ~�9t 2594t 46pw@�{�\sq ~�ΰ�q ~ q ~�9t 2595t 14pw@9K2�JBsq ~�ΰq ~ q ~�9t 2595t 15pw���:�㶚sq ~�ΰq ~ q ~�9t 2595t 43pw�ۘS��sq ~�ΰ�q ~ q ~�9t 2595t 49pw        sq ~�ΰ�q ~ q ~�9t 2596t 27pw@����tsq ~�ΰ�q ~ q ~�9t 2596t 68pw�����)�sq ~�ΰSq ~ q ~�9t 2597t 0pw@[���ssq ~�ΰ7q ~ q ~�9t 2597t 12pw��d��n�sq ~�ΰ�q ~ q ~�9t 2597t 22pw���)G��sq ~�ΰsq ~ q ~�9t 2597t 38pw��7�Ûsq ~�ΰ�q ~ q ~�9t 2597t 39pw?�/	߹sq ~�ΰ�q ~ q ~�9t 2597t 50pw        sq ~�ΰ�q ~ q ~�9t 2598t 12pw?�BX-b4sq ~�ΰWdq ~ q ~�9t 2598t 5pw        sq ~�ΰsq ~ q ~�9t 2599t 18pw?�<�O��sq ~�ΰ�q ~ q ~�9t 2599t 38pw        sq ~��W���q ~ q ~�9t 26t 0pw@7Xo9쬩sq ~��WŬq ~ q ~�9t 26t 12pw@C@yM��sq ~��WŬ�q ~ q ~�9t 26t 16pw?�"�>)�sq ~��Wů�q ~ q ~�9t 26t 22pw@@O�.S2sq ~��Wů�q ~ q ~�9t 26t 23pw        sq ~��Wų�q ~ q ~�9t 26t 32pw?��E��sq ~��Wŷ�q ~ q ~�9t 26t 46pw@�}���sq ~��W��q ~ q ~�9t 26t 5pw���txsq ~��Z��q ~ q ~�9t 260t 84pw@F�U�i�sq ~�ΰ�Xq ~ q ~�9t 2600t 14pw�����}sq ~�ΰ�wq ~ q ~�9t 2600t 15pw?����'�sq ~�ΰ�q ~ q ~�9t 2600t 72pw����u���sq ~�ΰ9�q ~ q ~�9t 2600t 8pw��bWrD�/sq ~�ΰ:q ~ q ~�9t 2600t 9pw?�y�u8u�sq ~�ΰ��q ~ q ~�9t 2601t 12pw?�4LcZ��sq ~�ΰ=fq ~ q ~�9t 2601t 6pw        sq ~�ΰ��q ~ q ~�9t 2602t 12pw?�4LcZ�usq ~�ΰ�q ~ q ~�9t 2602t 28pw        sq ~�ΰ�q ~ q ~�9t 2603t 84pw?�4LcZ�usq ~�ΰG�q ~ q ~�9t 2604t 0pw��I�1��sq ~�ΰ��q ~ q ~�9t 2604t 10pw        sq ~�ΰZq ~ q ~�9t 2604t 38pw@c��b$sq ~�ΰ�q ~ q ~�9t 2605t 12pw�����^sq ~�ΰ�q ~ q ~�9t 2605t 18pw?�.O��sq ~�ΰ:q ~ q ~�9t 2605t 39pw?��*��sq ~�ΰLKq ~ q ~�9t 2605t 5pw        sq ~�ΰ�q ~ q ~�9t 2606t 24pw��C���sq ~�ΰq ~ q ~�9t 2606t 31pw��k���sq ~�ΰq ~ q ~�9t 2606t 35pw���.YT|Nsq ~�ΰ�q ~ q ~�9t 2606t 52pw���.YT|Nsq ~�ΰ�q ~ q ~�9t 2606t 53pw��s2��Msq ~�ΰ�q ~ q ~�9t 2606t 54pw@��PF�sq ~�ΰ q ~ q ~�9t 2606t 67pw��½o%E�sq ~�ΰ`q ~ q ~�9t 2607t 24pw?�'���sq ~�ΰ�q ~ q ~�9t 2607t 31pw��4׌(��sq ~�ΰ@q ~ q ~�9t 2607t 35pw        sq ~�ΰ�q ~ q ~�9t 2607t 67pw�ݳ��oYsq ~�ΰ)�q ~ q ~�9t 2608t 84pw        sq ~�ΰ�q ~ q ~�9t 2609t 10pw        sq ~��Z��q ~ q ~�9t 261t 75pw        sq ~��Z��q ~ q ~�9t 261t 84pw@$      sq ~�ΰ�q ~ q ~�9t 2610t 84pw?���W-"sq ~�ΰ�q ~ q ~�9t 2611t 0pw����W�^sq ~�ΰqvq ~ q ~�9t 2611t 38pw?���>�`%sq ~�ΰt�q ~ q ~�9t 2611t 46pw        sq ~�ΰ��q ~ q ~�9t 2612t 84pw?��>�e sq ~�ΰt}q ~ q ~�9t 2613t 22pw?�p�9۪�sq ~�ΰ�q ~ q ~�9t 2613t 50pw        sq ~�ΰ�fq ~ q ~�9t 2613t 7pw�� 7®�0sq ~�ΰt�q ~ q ~�9t 2614t 14pw?�0W-�<Tsq ~�ΰt�q ~ q ~�9t 2614t 15pw��<�CPTsq ~�ΰx|q ~ q ~�9t 2615t 14pw?�Q�7���sq ~�ΰx�q ~ q ~�9t 2615t 15pw���r�h�sq ~�ΰ�bq ~ q ~�9t 2615t 41pw        sq ~�ΰ�q ~ q ~�9t 2615t 8pw��n��T@�sq ~�ΰ|=q ~ q ~�9t 2616t 14pw?�u�&�J�sq ~�ΰ|\q ~ q ~�9t 2616t 15pw��k��7%�sq ~�ΰ�q ~ q ~�9t 2616t 49pw        sq ~�ΰ��q ~ q ~�9t 2616t 72pw�Լ���sq ~�ΰ��q ~ q ~�9t 2616t 8pw?�.���sq ~�ΰ��q ~ q ~�9t 2616t 9pw��\|��_sq ~�ΰ�q ~ q ~�9t 2617t 12pw��O��o�sq ~�ΰ�zq ~ q ~�9t 2617t 18pw?��A�m�sq ~�ΰ��q ~ q ~�9t 2617t 37pw�zd�dYqsq ~�ΰ�q ~ q ~�9t 2617t 39pw        sq ~�ΰ�Gq ~ q ~�9t 2618t 50pw        sq ~�ΰ�q ~ q ~�9t 2618t 6pw?���O�sq ~�ΰ��q ~ q ~�9t 2619t 15pw?��a�Ȥsq ~�ΰ��q ~ q ~�9t 2619t 72pw        sq ~��Z� Iq ~ q ~�9t 262t 84pw@5oz�G�sq ~�ΰ�q ~ q ~�9t 2620t 14pw?�G.�sq ~�ΰ�5q ~ q ~�9t 2620t 15pw���&{u�sq ~�ΰ��q ~ q ~�9t 2620t 49pw        sq ~�ΰ�^q ~ q ~�9t 2620t 72pw�	�r���sq ~�ΰ"�q ~ q ~�9t 2620t 8pw��|�t�ڹsq ~�ΰ�[q ~ q ~�9t 2621t 10pw        sq ~�ΰ��q ~ q ~�9t 2621t 39pw?���+RJsq ~�ΰ�Wq ~ q ~�9t 2622t 48pw?޿��W[�sq ~�ΰ�q ~ q ~�9t 2623t 64pw?޿��W[�sq ~�ΰ��q ~ q ~�9t 2624t 61pw����.��sq ~�ΰ��q ~ q ~�9t 2624t 75pw        sq ~�ΰaq ~ q ~�9t 2624t 84pw?�WY�sq ~�ΰ�q ~ q ~�9t 2625t 16pw?�-���Csq ~�ΰ��q ~ q ~�9t 2625t 39pw        sq ~�ΰ�\q ~ q ~�9t 2625t 46pw?���?�sq ~�ΰ�q ~ q ~�9t 2626t 18pw�.���Vsq ~�ΰ�q ~ q ~�9t 2626t 22pw        sq ~�ΰ8�q ~ q ~�9t 2626t 6pw@n��l!_sq ~�ΰ�q ~ q ~�9t 2627t 55pw        sq ~�ΰ
�q ~ q ~�9t 2627t 73pw@@˜�	sq ~�ΰ��q ~ q ~�9t 2628t 24pw?�K�sq ~�ΰ@q ~ q ~�9t 2628t 67pw        sq ~�ΰ��q ~ q ~�9t 2629t 27pw?��G11��sq ~�ΰ(q ~ q ~�9t 2629t 60pw        sq ~��Z�$
q ~ q ~�9t 263t 84pw@F�U�i�sq ~�ΰR�q ~ q ~�9t 2630t 27pw@�c{Ĕsq ~�ΰ`�q ~ q ~�9t 2630t 60pw        sq ~�ΰR6q ~ q ~�9t 2631t 14pw���l�f�isq ~�ΰh~q ~ q ~�9t 2631t 72pw���,�D�sq ~�ΰ��q ~ q ~�9t 2631t 8pw��W�	v/sq ~�ΰV�q ~ q ~�9t 2632t 19pw@:��|sq ~�ΰ]Zq ~ q ~�9t 2632t 33pw�ƪ���gsq ~�ΰY�q ~ q ~�9t 2633t 14pw�����o�<sq ~�ΰY�q ~ q ~�9t 2633t 15pw@=�N�fsq ~�ΰd�q ~ q ~�9t 2633t 43pw����;��sq ~�ΰe�q ~ q ~�9t 2633t 49pw        sq ~�ΰa�q ~ q ~�9t 2634t 27pw?��O��sq ~�ΰa:q ~ q ~�9t 2635t 14pw?�F�ƴ�sq ~�ΰaYq ~ q ~�9t 2635t 15pw�r\��{QOsq ~�ΰmq ~ q ~�9t 2635t 49pw        sq ~�ΰw�q ~ q ~�9t 2635t 72pw��-�ݱB�sq ~�ΰ��q ~ q ~�9t 2635t 8pw?�^}??ksq ~�ΰ��q ~ q ~�9t 2635t 9pw����o�Tsq ~�ΰq ~ q ~�9t 2636t 82pw?��$l��sq ~�ΰ�Oq ~ q ~�9t 2637t 0pw?��$l��sq ~�ΰh�q ~ q ~�9t 2637t 16pw���IZR�>sq ~�ΰmq ~ q ~�9t 2637t 29pw        sq ~�ΰ��q ~ q ~�9t 2638t 73pw?����Ksq ~�ΰtq ~ q ~�9t 2639t 25pw?���sq ~�ΰ�q ~ q ~�9t 2639t 58pw        sq ~��Z�$)q ~ q ~�9t 264t 75pw        sq ~��Z�'�q ~ q ~�9t 264t 84pw@@�鹙�sq ~�ΰƕq ~ q ~�9t 2640t 24pw?�z���~�sq ~�ΰ��q ~ q ~�9t 2640t 71pw        sq ~�ΰƕq ~ q ~�9t 2641t 14pw�����sq ~�ΰƴq ~ q ~�9t 2641t 15pw?�W�#�?	sq ~�ΰ�sq ~ q ~�9t 2641t 49pw        sq ~�ΰ��q ~ q ~�9t 2641t 72pw���?���sq ~�ΰ q ~ q ~�9t 2641t 8pw��q�~~��sq ~�ΰ?q ~ q ~�9t 2641t 9pw?�Xf�W��sq ~�ΰ�q ~ q ~�9t 2642t 12pw?�s��-vsq ~�ΰβq ~ q ~�9t 2642t 29pw        sq ~�ΰ�q ~ q ~�9t 2643t 61pw        sq ~�ΰ�^q ~ q ~�9t 2643t 84pw?�s��-vsq ~�ΰ��q ~ q ~�9t 2644t 27pw?�����=�sq ~�ΰ�q ~ q ~�9t 2644t 68pw��X���sq ~�ΰՙq ~ q ~�9t 2645t 14pw��v����sq ~�ΰոq ~ q ~�9t 2645t 15pw�{%��I�$sq ~�ΰ�q ~ q ~�9t 2645t 41pw��HL[���sq ~�ΰ�q ~ q ~�9t 2645t 43pw���h���sq ~�ΰ�wq ~ q ~�9t 2645t 49pw        sq ~�ΰ��q ~ q ~�9t 2645t 72pw��/��f�sq ~�ΰ$q ~ q ~�9t 2645t 8pw@?)��6sq ~�ΰCq ~ q ~�9t 2645t 9pw���Ȧ�W�sq ~�ΰ�q ~ q ~�9t 2646t 31pw���2��ksq ~�ΰ� q ~ q ~�9t 2646t 52pw        sq ~�ΰ�|q ~ q ~�9t 2646t 67pw������ sq ~�ΰ�q ~ q ~�9t 2647t 14pw?��3{�s�sq ~�ΰ�cq ~ q ~�9t 2647t 72pw        sq ~�ΰ%�q ~ q ~�9t 2647t 8pw?��1��Vsq ~�ΰ�Dq ~ q ~�9t 2648t 61pw���9���Csq ~�ΰ�#q ~ q ~�9t 2648t 84pw?�;M�sq ~�ΰ,0q ~ q ~�9t 2649t 0pw��$�M�psq ~�ΰ�_q ~ q ~�9t 2649t 12pw��b�E�r�sq ~�ΰ,�q ~ q ~�9t 2649t 3pw?���QGsq ~�ΰ�q ~ q ~�9t 2649t 38pw        sq ~��Z�'�q ~ q ~�9t 265t 75pw        sq ~��Z�+�q ~ q ~�9t 265t 84pw@@�鹙�sq ~�ΰ~�q ~ q ~�9t 2650t 0pw��@�����sq ~�ΰ:�q ~ q ~�9t 2650t 22pw?�<�=adksq ~�ΰ?1q ~ q ~�9t 2650t 38pw?�;���k�sq ~�ΰE�q ~ q ~�9t 2650t 50pw        sq ~�ΰ:�q ~ q ~�9t 2651t 14pw��84��Busq ~�ΰ;q ~ q ~�9t 2651t 15pw�f���c77sq ~�ΰQ<q ~ q ~�9t 2651t 72pw��l�%sq ~�ΰ�q ~ q ~�9t 2651t 8pw@_OY�Xnsq ~�ΰ��q ~ q ~�9t 2651t 9pw�ןk@6E)sq ~�ΰM�q ~ q ~�9t 2652t 55pw        sq ~�ΰUq ~ q ~�9t 2652t 73pw@
��z��sq ~�ΰBWq ~ q ~�9t 2653t 13pw@��<�sq ~�ΰFuq ~ q ~�9t 2653t 26pw���	�1�sq ~�ΰJ6q ~ q ~�9t 2653t 36pw        sq ~�ΰM�q ~ q ~�9t 2653t 45pw��.����sq ~�ΰRq ~ q ~�9t 2653t 59pw��}��]sq ~�ΰ\�q ~ q ~�9t 2654t 73pw?��e�+sq ~�ΰI�q ~ q ~�9t 2655t 12pw��Z{=�csq ~�ΰN5q ~ q ~�9t 2655t 28pw        sq ~�ΰQ�q ~ q ~�9t 2656t 27pw        sq ~��Z�/Mq ~ q ~�9t 266t 84pw@@�鹙�sq ~��Z�/lq ~ q ~�9t 267t 75pw        sq ~��Z�3q ~ q ~�9t 267t 84pw@@�鹙�sq ~��Z�6�q ~ q ~�9t 268t 84pw@5oz�G�sq ~��Z�2�q ~ q ~�9t 269t 61pw        sq ~��Z�:�q ~ q ~�9t 269t 84pw@5oz�G�sq ~��Wų�q ~ q ~�9t 27t 24pw        sq ~��Wſq ~ q ~�9t 27t 54pw        sq ~��W��;q ~ q ~�9t 27t 67pw@$      sq ~��Z��&q ~ q ~�9t 270t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 271t 61pw        sq ~��Z���q ~ q ~�9t 271t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 272t 84pw@$      sq ~��Z���q ~ q ~�9t 273t 61pw        sq ~��Z��iq ~ q ~�9t 273t 84pw@@�鹙�sq ~��Z��Kq ~ q ~�9t 274t 61pw        sq ~��Z��*q ~ q ~�9t 274t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 275t 61pw        sq ~��Z���q ~ q ~�9t 275t 84pw@$      sq ~��Z���q ~ q ~�9t 276t 61pw        sq ~��Z���q ~ q ~�9t 276t 84pw@5oz�G�sq ~��Z��mq ~ q ~�9t 277t 84pw@@�鹙�sq ~��Z��Oq ~ q ~�9t 278t 61pw        sq ~��Z��.q ~ q ~�9t 278t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 279t 84pw@@�鹙�sq ~��Wŷ�q ~ q ~�9t 28t 25pw        sq ~��Wź�q ~ q ~�9t 28t 30pw@5oz�G�sq ~��W��;q ~ q ~�9t 28t 57pw@5oz�G�sq ~��Z���q ~ q ~�9t 280t 75pw        sq ~��Z��q ~ q ~�9t 280t 84pw@$      sq ~��Z��gq ~ q ~�9t 281t 61pw        sq ~��Z�Fq ~ q ~�9t 281t 84pw@@�鹙�sq ~��Z�eq ~ q ~�9t 282t 75pw        sq ~��Z�	q ~ q ~�9t 282t 84pw@5oz�G�sq ~��Z�	&q ~ q ~�9t 283t 75pw        sq ~��Z��q ~ q ~�9t 283t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 284t 75pw        sq ~��Z��q ~ q ~�9t 284t 84pw@F�U�i�sq ~��Z�kq ~ q ~�9t 285t 61pw        sq ~��Z�Jq ~ q ~�9t 285t 84pw@$      sq ~��Z�,q ~ q ~�9t 286t 61pw        sq ~��Z�q ~ q ~�9t 286t 84pw@$      sq ~��Z��q ~ q ~�9t 287t 61pw        sq ~��Z��q ~ q ~�9t 287t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 288t 61pw        sq ~��Z��q ~ q ~�9t 288t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 289t 75pw        sq ~��Z�#Nq ~ q ~�9t 289t 84pw@$      sq ~��WŻ�q ~ q ~�9t 29t 27pw        sq ~��W���q ~ q ~�9t 29t 68pw@+�Ք��sq ~��Z�rBq ~ q ~�9t 290t 75pw        sq ~��Z�u�q ~ q ~�9t 290t 84pw@5oz�G�sq ~��Z�vq ~ q ~�9t 291t 75pw        sq ~��Z�y�q ~ q ~�9t 291t 84pw@5oz�G�sq ~��Z�}fq ~ q ~�9t 292t 84pw@@�鹙�sq ~��Z�yHq ~ q ~�9t 293t 61pw        sq ~��Z��'q ~ q ~�9t 293t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 294t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 295t 84pw@M]��%��sq ~��Z��jq ~ q ~�9t 296t 84pw@@�鹙�sq ~��Z��Lq ~ q ~�9t 297t 61pw        sq ~��Z��+q ~ q ~�9t 297t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 298t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 299t 84pw@5oz�G�sq ~��W���q ~ q ~�9t 3t 21pw@$      sq ~��W��q ~ q ~�9t 3t 26pw        sq ~��W�.�q ~ q ~�9t 3t 4pw        sq ~��W�	�q ~ q ~�9t 30t 12pw?����v�sq ~��W�nq ~ q ~�9t 30t 28pw        sq ~��W�R_q ~ q ~�9t 30t 5pw@4p$�@�sq ~��Z�vq ~ q ~�9t 300t 84pw@@�鹙�sq ~��Z�q�q ~ q ~�9t 301t 61pw        sq ~��Z�y�q ~ q ~�9t 301t 84pw@5oz�G�sq ~��Z�}�q ~ q ~�9t 302t 84pw@$      sq ~��Z�yrq ~ q ~�9t 303t 61pw        sq ~��Z��Qq ~ q ~�9t 303t 84pw@F�U�i�sq ~��Z��q ~ q ~�9t 304t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 305t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 306t 84pw@F�U�i�sq ~��Z��Uq ~ q ~�9t 307t 84pw@F�U�i�sq ~��Z��7q ~ q ~�9t 308t 61pw        sq ~��Z��q ~ q ~�9t 308t 84pw@@�鹙�sq ~��Z��5q ~ q ~�9t 309t 75pw        sq ~��Z���q ~ q ~�9t 309t 84pw@@�鹙�sq ~��W�q ~ q ~�9t 31t 31pw        sq ~��W��q ~ q ~�9t 31t 35pw        sq ~��W�!q ~ q ~�9t 31t 67pw@$�ε��sq ~��Z���q ~ q ~�9t 310t 75pw        sq ~��Z��mq ~ q ~�9t 310t 84pw@5oz�G�sq ~��Z��Oq ~ q ~�9t 311t 61pw        sq ~��Z��.q ~ q ~�9t 311t 84pw@5oz�G�sq ~��Z��Mq ~ q ~�9t 312t 75pw        sq ~��Z���q ~ q ~�9t 312t 84pw@$      sq ~��Z���q ~ q ~�9t 313t 84pw@#�i����sq ~��Z���q ~ q ~�9t 314t 75pw        sq ~��Z��qq ~ q ~�9t 314t 84pw@5oz�G�sq ~��Z��2q ~ q ~�9t 315t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 316t 61pw        sq ~��Z� �q ~ q ~�9t 316t 84pw@$      sq ~��Z���q ~ q ~�9t 317t 61pw        sq ~��Z��q ~ q ~�9t 317t 84pw@5oz�G�sq ~��Z� �q ~ q ~�9t 318t 61pw        sq ~��Z�uq ~ q ~�9t 318t 84pw@@�鹙�sq ~��Z�Wq ~ q ~�9t 319t 61pw�1+���ksq ~��Z�6q ~ q ~�9t 319t 84pw@)�A>hA	sq ~��W�Y�q ~ q ~�9t 32t 2pw        sq ~��W�q ~ q ~�9t 32t 21pw@$      sq ~��W�Y�q ~ q ~�9t 32t 4pw@$      sq ~��W��q ~ q ~�9t 32t 44pw        sq ~��W�!Rq ~ q ~�9t 32t 59pw@$      sq ~��Z�[*q ~ q ~�9t 320t 75pw        sq ~��Z�^�q ~ q ~�9t 320t 84pw@5oz�G�sq ~��Z�^�q ~ q ~�9t 321t 75pw        sq ~��Z�b�q ~ q ~�9t 321t 84pw@F�U�i�sq ~��Z�fNq ~ q ~�9t 322t 84pw@5oz�G�sq ~��Z�b0q ~ q ~�9t 323t 61pw        sq ~��Z�jq ~ q ~�9t 323t 84pw@5oz�G�sq ~��Z�e�q ~ q ~�9t 324t 61pw        sq ~��Z�m�q ~ q ~�9t 324t 84pw@@�鹙�sq ~��Z�q�q ~ q ~�9t 325t 84pw@@�鹙�sq ~��Z�uRq ~ q ~�9t 326t 84pw@$      sq ~��Z�uqq ~ q ~�9t 327t 75pw        sq ~��Z�yq ~ q ~�9t 327t 84pw@5oz�G�sq ~��Z�t�q ~ q ~�9t 328t 61pw        sq ~��Z�|�q ~ q ~�9t 328t 84pw@$      sq ~��Z�|�q ~ q ~�9t 329t 75pw        sq ~��Z���q ~ q ~�9t 329t 84pw@$      sq ~��W�q ~ q ~�9t 33t 19pw@5oz�G�sq ~��W��q ~ q ~�9t 33t 33pw        sq ~��W�(q ~ q ~�9t 33t 63pw        sq ~��Z�ωq ~ q ~�9t 330t 75pw        sq ~��Z��+q ~ q ~�9t 330t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 331t 84pw@$      sq ~��Z�ڭq ~ q ~�9t 332t 84pw@5oz�G�sq ~��Z��nq ~ q ~�9t 333t 84pw@@�鹙�sq ~��Z��/q ~ q ~�9t 334t 84pw@5oz�G�sq ~��Z��Nq ~ q ~�9t 335t 75pw        sq ~��Z���q ~ q ~�9t 335t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 336t 84pw@@�鹙�sq ~��Z��rq ~ q ~�9t 337t 84pw@$      sq ~��Z��3q ~ q ~�9t 338t 84pw@$      sq ~��Z��Rq ~ q ~�9t 339t 75pw        sq ~��Z���q ~ q ~�9t 339t 84pw@5oz�G�sq ~��W�aq ~ q ~�9t 34t 2pw@$J_X6��sq ~��W��q ~ q ~�9t 34t 21pw?��*rK@sq ~��W� �q ~ q ~�9t 34t 34pw        sq ~��Z�G�q ~ q ~�9t 340t 84pw@5oz�G�sq ~��Z�KKq ~ q ~�9t 341t 84pw@$      sq ~��Z�G-q ~ q ~�9t 342t 61pw        sq ~��Z�Oq ~ q ~�9t 342t 84pw@5oz�G�sq ~��Z�R�q ~ q ~�9t 343t 84pw@@�鹙�sq ~��Z�N�q ~ q ~�9t 344t 61pw        sq ~��Z�V�q ~ q ~�9t 344t 84pw@$      sq ~��Z�ZOq ~ q ~�9t 345t 84pw@5oz�G�sq ~��Z�V1q ~ q ~�9t 346t 61pw        sq ~��Z�^q ~ q ~�9t 346t 84pw@@�鹙�sq ~��Z�^/q ~ q ~�9t 347t 75pw        sq ~��Z�a�q ~ q ~�9t 347t 84pw@$      sq ~��Z�a�q ~ q ~�9t 348t 75pw        sq ~��Z�e�q ~ q ~�9t 348t 84pw@@�鹙�sq ~��Z�atq ~ q ~�9t 349t 61pw        sq ~��Z�iSq ~ q ~�9t 349t 84pw@$      sq ~��W��q ~ q ~�9t 35t 13pw@%�1��Msq ~��W�$�q ~ q ~�9t 35t 36pw        sq ~��Z��Gq ~ q ~�9t 350t 75pw        sq ~��Z���q ~ q ~�9t 350t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 351t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 352t 75pw        sq ~��Z��kq ~ q ~�9t 352t 84pw@$      sq ~��Z��Mq ~ q ~�9t 353t 61pw        sq ~��Z��,q ~ q ~�9t 353t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 354t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 355t 75pw        sq ~��Z�ήq ~ q ~�9t 355t 84pw@F�U�i�sq ~��Z��oq ~ q ~�9t 356t 84pw@F�U�i�sq ~��Z�Ҏq ~ q ~�9t 357t 75pw        sq ~��Z��0q ~ q ~�9t 357t 84pw@5oz�G�sq ~��Z��Oq ~ q ~�9t 358t 75pw        sq ~��Z���q ~ q ~�9t 358t 84pw@$      sq ~��Z���q ~ q ~�9t 359t 61pw        sq ~��Z�ݲq ~ q ~�9t 359t 84pw@5oz�G�sq ~��W�hJq ~ q ~�9t 36t 0pw����j�%�sq ~��W� yq ~ q ~�9t 36t 12pw�������sq ~��W� �q ~ q ~�9t 36t 16pw��5�޴�[sq ~��W�$:q ~ q ~�9t 36t 22pw@#{��sq ~��W�$�q ~ q ~�9t 36t 28pw��o1�p(�sq ~��W�'�q ~ q ~�9t 36t 32pw��H��H�sq ~��W�,8q ~ q ~�9t 36t 46pw��L�Y`�nsq ~��W�h�q ~ q ~�9t 36t 5pw        sq ~��Z�,�q ~ q ~�9t 360t 75pw        sq ~��Z�0Hq ~ q ~�9t 360t 84pw@@�鹙�sq ~��Z�4	q ~ q ~�9t 361t 84pw@@�鹙�sq ~��Z�7�q ~ q ~�9t 362t 84pw@@�鹙�sq ~��Z�;�q ~ q ~�9t 363t 84pw@@�鹙�sq ~��Z�7mq ~ q ~�9t 364t 61pw        sq ~��Z�?Lq ~ q ~�9t 364t 84pw@@�鹙�sq ~��Z�Cq ~ q ~�9t 365t 84pw@$      sq ~��Z�F�q ~ q ~�9t 366t 84pw@F�U�i�sq ~��Z�B�q ~ q ~�9t 367t 61pw        sq ~��Z�J�q ~ q ~�9t 367t 84pw@5oz�G�sq ~��Z�Fqq ~ q ~�9t 368t 61pw        sq ~��Z�NPq ~ q ~�9t 368t 84pw@5oz�G�sq ~��Z�J2q ~ q ~�9t 369t 61pw        sq ~��Z�Rq ~ q ~�9t 369t 84pw@5oz�G�sq ~��W�/?q ~ q ~�9t 37t 40pw        sq ~��W�3�q ~ q ~�9t 37t 58pw@$      sq ~��W�7�q ~ q ~�9t 37t 69pw@$      sq ~��Z���q ~ q ~�9t 370t 61pw        sq ~��Z���q ~ q ~�9t 370t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 371t 61pw        sq ~��Z��hq ~ q ~�9t 371t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 372t 75pw        sq ~��Z��)q ~ q ~�9t 372t 84pw@@�鹙�sq ~��Z��Hq ~ q ~�9t 373t 75pw        sq ~��Z���q ~ q ~�9t 373t 84pw@F�U�i�sq ~��Z��	q ~ q ~�9t 374t 75pw        sq ~��Z���q ~ q ~�9t 374t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 375t 61pw        sq ~��Z��lq ~ q ~�9t 375t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 376t 75pw        sq ~��Z��-q ~ q ~�9t 376t 84pw@$      sq ~��Z��q ~ q ~�9t 377t 61pw        sq ~��Z���q ~ q ~�9t 377t 84pw@$F�\#=�sq ~��Z�¯q ~ q ~�9t 378t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 379t 75pw        sq ~��Z��pq ~ q ~�9t 379t 84pw@$      sq ~��W�07q ~ q ~�9t 38t 38pw@5oz�G�sq ~��W�p�q ~ q ~�9t 38t 6pw        sq ~��Z�q ~ q ~�9t 380t 84pw@@�鹙�sq ~��Z�%q ~ q ~�9t 381t 75pw        sq ~��Z��q ~ q ~�9t 381t 84pw@$      sq ~��Z��q ~ q ~�9t 382t 61pw        sq ~��Z� �q ~ q ~�9t 382t 84pw@@�鹙�sq ~��Z�$Iq ~ q ~�9t 383t 84pw@$      sq ~��Z� +q ~ q ~�9t 384t 61pw        sq ~��Z�(
q ~ q ~�9t 384t 84pw@@�鹙�sq ~��Z�+�q ~ q ~�9t 385t 84pw@$      sq ~��Z�'�q ~ q ~�9t 386t 61pw        sq ~��Z�/�q ~ q ~�9t 386t 84pw@@�鹙�sq ~��Z�3Mq ~ q ~�9t 387t 84pw@$      sq ~��Z�//q ~ q ~�9t 388t 61pw        sq ~��Z�7q ~ q ~�9t 388t 84pw@@�鹙�sq ~��Z�:�q ~ q ~�9t 389t 84pw@F�U�i�sq ~��W�3q ~ q ~�9t 39t 31pw        sq ~��W�3�q ~ q ~�9t 39t 35pw@5oz�G�sq ~��W�:�q ~ q ~�9t 39t 52pw@5oz�G�sq ~��W�B#q ~ q ~�9t 39t 71pw        sq ~��Z���q ~ q ~�9t 390t 61pw        sq ~��Z��eq ~ q ~�9t 390t 84pw@$��ɶ�sq ~��Z��&q ~ q ~�9t 391t 84pw@5oz�G�sq ~��Z��Eq ~ q ~�9t 392t 75pw        sq ~��Z���q ~ q ~�9t 392t 84pw@$      sq ~��Z���q ~ q ~�9t 393t 84pw@$      sq ~��Z���q ~ q ~�9t 394t 75pw        sq ~��Z��iq ~ q ~�9t 394t 84pw@$      sq ~��Z��Kq ~ q ~�9t 395t 61pw        sq ~��Z��*q ~ q ~�9t 395t 84pw@5oz�G�sq ~��Z��Iq ~ q ~�9t 396t 75pw        sq ~��Z���q ~ q ~�9t 396t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 397t 61pw        sq ~��Z���q ~ q ~�9t 397t 84pw@$      sq ~��Z���q ~ q ~�9t 398t 61pw        sq ~��Z��mq ~ q ~�9t 398t 84pw@5oz�G�sq ~��Z��Oq ~ q ~�9t 399t 61pw        sq ~��Z��.q ~ q ~�9t 399t 84pw@5oz�G�sq ~��W�1�q ~ q ~�9t 4t 0pw���"6sq ~��W��
q ~ q ~�9t 4t 12pw��;}��sq ~��W���q ~ q ~�9t 4t 22pw@��-gD%sq ~��W��q ~ q ~�9t 4t 28pw@,衘�~�sq ~��W�28q ~ q ~�9t 4t 3pw@ E���[sq ~��W��q ~ q ~�9t 4t 32pw@$^�����sq ~��W�2vq ~ q ~�9t 4t 5pw        sq ~��W���q ~ q ~�9t 4t 50pw@%�����$sq ~��W�2�q ~ q ~�9t 4t 6pw?�k�#��'sq ~��W�~�q ~ q ~�9t 40t 14pw@)��bp��sq ~��WƉvq ~ q ~�9t 40t 41pw        sq ~��WƔ�q ~ q ~�9t 40t 72pw�a��-��sq ~��Z���q ~ q ~�9t 400t 75pw        sq ~��Z���q ~ q ~�9t 400t 84pw@5oz�G�sq ~��Z��Pq ~ q ~�9t 401t 84pw@5x�E�sq ~��Z��q ~ q ~�9t 402t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 403t 61pw        sq ~��Z���q ~ q ~�9t 403t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 404t 75pw        sq ~��Z���q ~ q ~�9t 404t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 405t 75pw        sq ~��Z��Tq ~ q ~�9t 405t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 406t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 407t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 408t 75pw        sq ~��Z���q ~ q ~�9t 408t 84pw@@�鹙�sq ~��Z��Xq ~ q ~�9t 409t 84pw@5oz�G�sq ~��WƂ2q ~ q ~�9t 41t 13pw���=h��
sq ~��Wƅ�q ~ q ~�9t 41t 21pw@$      sq ~��WƆPq ~ q ~�9t 41t 26pw� 9�! �sq ~��W��`q ~ q ~�9t 41t 4pw@$����sq ~��WƍVq ~ q ~�9t 41t 42pw        sq ~��Wƍ�q ~ q ~�9t 41t 45pw� ���" �sq ~��WƑ�q ~ q ~�9t 41t 59pw@%�iƲsq ~��Z��q ~ q ~�9t 410t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 411t 84pw@5oz�G�sq ~��Z�	pq ~ q ~�9t 412t 84pw@@�鹙�sq ~��Z�1q ~ q ~�9t 413t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 414t 84pw@$      sq ~��Z��q ~ q ~�9t 415t 61pw        sq ~��Z��q ~ q ~�9t 415t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 416t 61pw        sq ~��Z�tq ~ q ~�9t 416t 84pw@5oz�G�sq ~��Z�Vq ~ q ~�9t 417t 61pw        sq ~��Z�5q ~ q ~�9t 417t 84pw@$      sq ~��Z�q ~ q ~�9t 418t 61pw        sq ~��Z��q ~ q ~�9t 418t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 419t 61pw        sq ~��Z�#�q ~ q ~�9t 419t 84pw@F�U�i�sq ~��WƆ1q ~ q ~�9t 42t 15pw@'3k�wV�sq ~��WƑ6q ~ q ~�9t 42t 43pw        sq ~��Z�r�q ~ q ~�9t 420t 75pw        sq ~��Z�vMq ~ q ~�9t 420t 84pw@5oz�G�sq ~��Z�zq ~ q ~�9t 421t 84pw@%�k԰�sq ~��Z�}�q ~ q ~�9t 422t 84pw@5oz�G�sq ~��Z�}�q ~ q ~�9t 423t 75pw        sq ~��Z���q ~ q ~�9t 423t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 424t 75pw        sq ~��Z��Qq ~ q ~�9t 424t 84pw@$      sq ~��Z��3q ~ q ~�9t 425t 61pw        sq ~��Z��q ~ q ~�9t 425t 84pw@%���}B�sq ~��Z���q ~ q ~�9t 426t 61pw        sq ~��Z���q ~ q ~�9t 426t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 427t 75pw        sq ~��Z���q ~ q ~�9t 427t 84pw@5oz�G�sq ~��Z��Uq ~ q ~�9t 428t 84pw@F�U�i�sq ~��Z��7q ~ q ~�9t 429t 61pw        sq ~��Z��q ~ q ~�9t 429t 84pw@@�鹙�sq ~��W��fq ~ q ~�9t 43t 0pw��,��:��sq ~��WƉ�q ~ q ~�9t 43t 12pw@8,�� O�sq ~��WƍVq ~ q ~�9t 43t 22pw@&�� ��ysq ~��W���q ~ q ~�9t 43t 3pw��I�1��sq ~��WƑ�q ~ q ~�9t 43t 38pw        sq ~��WƑ�q ~ q ~�9t 43t 39pw?��*�}sq ~��W��?q ~ q ~�9t 43t 7pw@%Y����zsq ~��Z���q ~ q ~�9t 430t 61pw        sq ~��Z��q ~ q ~�9t 430t 84pw@5oz�G�sq ~��Z��mq ~ q ~�9t 431t 84pw@$      sq ~��Z��q ~ q ~�9t 432t 75pw        sq ~��Z��.q ~ q ~�9t 432t 84pw@5oz�G�sq ~��Z��Mq ~ q ~�9t 433t 75pw        sq ~��Z���q ~ q ~�9t 433t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 434t 84pw@5oz�G�sq ~��Z��qq ~ q ~�9t 435t 84pw@5oz�G�sq ~��Z�2q ~ q ~�9t 436t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 437t 61pw        sq ~��Z��q ~ q ~�9t 437t 84pw@@�鹙�sq ~��Z� �q ~ q ~�9t 438t 61pw        sq ~��Z��q ~ q ~�9t 438t 84pw@@�鹙�sq ~��Z�uq ~ q ~�9t 439t 84pw@@�鹙�sq ~��WƘzq ~ q ~�9t 44t 41pw        sq ~��Wƙrq ~ q ~�9t 44t 49pw@5oz�G�sq ~��Z�W,q ~ q ~�9t 440t 61pw        sq ~��Z�_q ~ q ~�9t 440t 84pw@5oz�G�sq ~��Z�Z�q ~ q ~�9t 441t 61pw        sq ~��Z�b�q ~ q ~�9t 441t 84pw@5oz�G�sq ~��Z�b�q ~ q ~�9t 442t 75pw        sq ~��Z�f�q ~ q ~�9t 442t 84pw@@�鹙�sq ~��Z�boq ~ q ~�9t 443t 61pw        sq ~��Z�jNq ~ q ~�9t 443t 84pw@5oz�G�sq ~��Z�f0q ~ q ~�9t 444t 61pw        sq ~��Z�nq ~ q ~�9t 444t 84pw@$      sq ~��Z�n.q ~ q ~�9t 445t 75pw        sq ~��Z�q�q ~ q ~�9t 445t 84pw@5oz�G�sq ~��Z�u�q ~ q ~�9t 446t 84pw@5oz�G�sq ~��Z�u�q ~ q ~�9t 447t 75pw        sq ~��Z�yRq ~ q ~�9t 447t 84pw@5oz�G�sq ~��Z�}q ~ q ~�9t 448t 84pw@@�鹙�sq ~��Z�}2q ~ q ~�9t 449t 75pw        sq ~��Z���q ~ q ~�9t 449t 84pw@#3^-��sq ~��WƑ�q ~ q ~�9t 45t 19pw?�5�?�Y�sq ~��WƘ�q ~ q ~�9t 45t 33pw��M�#sq ~��Wƣ�q ~ q ~�9t 45t 63pw@%���t�sq ~��WƤ9q ~ q ~�9t 45t 65pw@%.���2sq ~��Z�ˋq ~ q ~�9t 450t 61pw        sq ~��Z��jq ~ q ~�9t 450t 84pw@$      sq ~��Z��+q ~ q ~�9t 451t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 452t 84pw@$      sq ~��Z���q ~ q ~�9t 453t 61pw        sq ~��Z�ޭq ~ q ~�9t 453t 84pw@$      sq ~��Z��nq ~ q ~�9t 454t 84pw@F�U�i�sq ~��Z��Pq ~ q ~�9t 455t 61pw        sq ~��Z��/q ~ q ~�9t 455t 84pw@@�鹙�sq ~��Z��Nq ~ q ~�9t 456t 75pw        sq ~��Z���q ~ q ~�9t 456t 84pw@"5w�*sq ~��Z��q ~ q ~�9t 457t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 458t 75pw        sq ~��Z��rq ~ q ~�9t 458t 84pw@@�鹙�sq ~��Z��3q ~ q ~�9t 459t 84pw@F�U�i�sq ~��WƘzq ~ q ~�9t 46t 21pw@0�z�:�wsq ~��Wƙq ~ q ~�9t 46t 26pw@&�Bk��sq ~��WƜ�q ~ q ~�9t 46t 34pw@$      sq ~��WƜ�q ~ q ~�9t 46t 36pw@���ssq ~��W��%q ~ q ~�9t 46t 4pw���o�*��sq ~��WƠYq ~ q ~�9t 46t 44pw@#��!��sq ~��WƤ�q ~ q ~�9t 46t 59pw���ꚻ�sq ~��Z�D'q ~ q ~�9t 460t 75pw        sq ~��Z�G�q ~ q ~�9t 460t 84pw@5oz�G�sq ~��Z�C�q ~ q ~�9t 461t 61pw        sq ~��Z�K�q ~ q ~�9t 461t 84pw@5oz�G�sq ~��Z�K�q ~ q ~�9t 462t 75pw        sq ~��Z�OKq ~ q ~�9t 462t 84pw@@�鹙�sq ~��Z�Ojq ~ q ~�9t 463t 75pw        sq ~��Z�Sq ~ q ~�9t 463t 84pw@5oz�G�sq ~��Z�N�q ~ q ~�9t 464t 61pw        sq ~��Z�V�q ~ q ~�9t 464t 84pw@5oz�G�sq ~��Z�V�q ~ q ~�9t 465t 75pw        sq ~��Z�Z�q ~ q ~�9t 465t 84pw@5oz�G�sq ~��Z�Vpq ~ q ~�9t 466t 61pw        sq ~��Z�^Oq ~ q ~�9t 466t 84pw@F�U�i�sq ~��Z�^nq ~ q ~�9t 467t 75pw        sq ~��Z�bq ~ q ~�9t 467t 84pw@@�鹙�sq ~��Z�]�q ~ q ~�9t 468t 61pw        sq ~��Z�e�q ~ q ~�9t 468t 84pw@@�鹙�sq ~��Z�a�q ~ q ~�9t 469t 61pw        sq ~��Z�i�q ~ q ~�9t 469t 84pw@5oz�G�sq ~��WƘ�q ~ q ~�9t 47t 13pw��HI�h�sq ~��WƜ;q ~ q ~�9t 47t 21pw@$      sq ~��WƜ�q ~ q ~�9t 47t 26pw�����<��sq ~��WƤ9q ~ q ~�9t 47t 45pw��ruo��sq ~��Z���q ~ q ~�9t 470t 75pw        sq ~��Z��(q ~ q ~�9t 470t 84pw@5oz�G�sq ~��Z��Gq ~ q ~�9t 471t 75pw        sq ~��Z���q ~ q ~�9t 471t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 472t 61pw        sq ~��Z�êq ~ q ~�9t 472t 84pw@$      sq ~��Z���q ~ q ~�9t 473t 75pw        sq ~��Z��kq ~ q ~�9t 473t 84pw@@�鹙�sq ~��Z�Ǌq ~ q ~�9t 474t 75pw        sq ~��Z��,q ~ q ~�9t 474t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 475t 61pw        sq ~��Z���q ~ q ~�9t 475t 84pw@5oz�G�sq ~��Z�Үq ~ q ~�9t 476t 84pw@$      sq ~��Z�ΐq ~ q ~�9t 477t 61pw        sq ~��Z��oq ~ q ~�9t 477t 84pw@$      sq ~��Z��0q ~ q ~�9t 478t 84pw@$      sq ~��Z��Oq ~ q ~�9t 479t 75pw        sq ~��Z���q ~ q ~�9t 479t 84pw@5oz�G�sq ~��WƜZq ~ q ~�9t 48t 12pw��1Jesq ~��WƜ�q ~ q ~�9t 48t 16pw?���E�sq ~��WƠ�q ~ q ~�9t 48t 28pw?�ˎ��sq ~��W��q ~ q ~�9t 48t 3pw@&�C"{i�sq ~��Wƣ�q ~ q ~�9t 48t 32pw?�rLA���sq ~��Wƨq ~ q ~�9t 48t 46pw?�1� �),sq ~��W���q ~ q ~�9t 48t 5pw        sq ~��Z�(�q ~ q ~�9t 480t 61pw        sq ~��Z�0�q ~ q ~�9t 480t 84pw@5oz�G�sq ~��Z�4Hq ~ q ~�9t 481t 84pw@$      sq ~��Z�0*q ~ q ~�9t 482t 61pw        sq ~��Z�8	q ~ q ~�9t 482t 84pw@F�U�i�sq ~��Z�8(q ~ q ~�9t 483t 75pw        sq ~��Z�;�q ~ q ~�9t 483t 84pw@$      sq ~��Z�;�q ~ q ~�9t 484t 75pw        sq ~��Z�?�q ~ q ~�9t 484t 84pw@$      sq ~��Z�;mq ~ q ~�9t 485t 61pw        sq ~��Z�CLq ~ q ~�9t 485t 84pw@5oz�G�sq ~��Z�Gq ~ q ~�9t 486t 84pw@5oz�G�sq ~��Z�J�q ~ q ~�9t 487t 84pw@$      sq ~��Z�J�q ~ q ~�9t 488t 75pw        sq ~��Z�N�q ~ q ~�9t 488t 84pw@$      sq ~��Z�RPq ~ q ~�9t 489t 84pw@@�鹙�sq ~��W��q ~ q ~�9t 49t 1pw@&��+Asq ~��WƳ\q ~ q ~�9t 49t 66pw@$      sq ~��Z��Dq ~ q ~�9t 490t 75pw        sq ~��Z���q ~ q ~�9t 490t 84pw@#���*�sq ~��Z���q ~ q ~�9t 491t 61pw        sq ~��Z���q ~ q ~�9t 491t 84pw@@�鹙�sq ~��Z��hq ~ q ~�9t 492t 84pw@$      sq ~��Z��Jq ~ q ~�9t 493t 61pw        sq ~��Z��)q ~ q ~�9t 493t 84pw@F�U�i�sq ~��Z��q ~ q ~�9t 494t 61pw        sq ~��Z���q ~ q ~�9t 494t 84pw@@�鹙�sq ~��Z��	q ~ q ~�9t 495t 75pw        sq ~��Z���q ~ q ~�9t 495t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 496t 61pw        sq ~��Z��lq ~ q ~�9t 496t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 497t 75pw        sq ~��Z��-q ~ q ~�9t 497t 84pw@@�鹙�sq ~��Z��Lq ~ q ~�9t 498t 75pw        sq ~��Z���q ~ q ~�9t 498t 84pw@@�鹙�sq ~��Z�Ưq ~ q ~�9t 499t 84pw@5oz�G�sq ~��W��Gq ~ q ~�9t 5t 16pw?л[�`isq ~��W��q ~ q ~�9t 5t 23pw@$      sq ~��W��Fq ~ q ~�9t 5t 28pw���s2m}sq ~��W��Mq ~ q ~�9t 5t 32pw���/�{�sq ~��W��q ~ q ~�9t 5t 38pw?�K�sq ~��W���q ~ q ~�9t 5t 46pw?�5^�MRsq ~��W�6uq ~ q ~�9t 5t 7pw        sq ~��W���q ~ q ~�9t 50t 24pw�h����Wsq ~��W��q ~ q ~�9t 50t 53pw        sq ~��W�q ~ q ~�9t 50t 67pw@#�0�D7jsq ~��W�	q ~ q ~�9t 50t 71pw@$      sq ~��Z��nq ~ q ~�9t 500t 75pw        sq ~��Z��q ~ q ~�9t 500t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 501t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 502t 61pw        sq ~��Z���q ~ q ~�9t 502t 84pw@5oz�G�sq ~��Z��tq ~ q ~�9t 503t 61pw        sq ~��Z��Sq ~ q ~�9t 503t 84pw@@�鹙�sq ~��Z��rq ~ q ~�9t 504t 75pw        sq ~��Z��q ~ q ~�9t 504t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 505t 61pw        sq ~��Z���q ~ q ~�9t 505t 84pw@$      sq ~��Z���q ~ q ~�9t 506t 61pw        sq ~��Z���q ~ q ~�9t 506t 84pw@@�鹙�sq ~��Z��Wq ~ q ~�9t 507t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 508t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 509t 61pw        sq ~��Z���q ~ q ~�9t 509t 84pw@$      sq ~��W���q ~ q ~�9t 51t 14pw@0��,�%Rsq ~��W���q ~ q ~�9t 51t 20pw        sq ~��Z��q ~ q ~�9t 510t 61pw        sq ~��Z�oq ~ q ~�9t 510t 84pw@$      sq ~��Z�0q ~ q ~�9t 511t 84pw@@�鹙�sq ~��Z�Oq ~ q ~�9t 512t 75pw        sq ~��Z� �q ~ q ~�9t 512t 84pw@@�鹙�sq ~��Z�$�q ~ q ~�9t 513t 84pw@5oz�G�sq ~��Z� �q ~ q ~�9t 514t 61pw        sq ~��Z�(sq ~ q ~�9t 514t 84pw@@�鹙�sq ~��Z�,4q ~ q ~�9t 515t 84pw@@�鹙�sq ~��Z�/�q ~ q ~�9t 516t 84pw@5oz�G�sq ~��Z�3�q ~ q ~�9t 517t 84pw@$      sq ~��Z�3�q ~ q ~�9t 518t 75pw        sq ~��Z�7wq ~ q ~�9t 518t 84pw@5oz�G�sq ~��Z�;8q ~ q ~�9t 519t 84pw@5oz�G�sq ~��W�0q ~ q ~�9t 52t 48pw@5oz�G�sq ~��Z���q ~ q ~�9t 520t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 521t 61pw        sq ~��Z���q ~ q ~�9t 521t 84pw@@�鹙�sq ~��Z��Pq ~ q ~�9t 522t 84pw@5oz�G�sq ~��Z��oq ~ q ~�9t 523t 75pw        sq ~��Z��q ~ q ~�9t 523t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 524t 84pw@$&L��@sq ~��Z���q ~ q ~�9t 525t 75pw        sq ~��Z���q ~ q ~�9t 525t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 526t 75pw        sq ~��Z��Tq ~ q ~�9t 526t 84pw@5oz�G�sq ~��Z��6q ~ q ~�9t 527t 61pw        sq ~��Z��q ~ q ~�9t 527t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 528t 61pw        sq ~��Z���q ~ q ~�9t 528t 84pw@$      sq ~��Z���q ~ q ~�9t 529t 84pw@F�U�i�sq ~��W��q ~ q ~�9t 53t 24pw����d�sq ~��W�Wq ~ q ~�9t 53t 31pw@&k�sq ~��Z��Nq ~ q ~�9t 530t 61pw        sq ~��Z�-q ~ q ~�9t 530t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 531t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 532t 61pw        sq ~��Z�	�q ~ q ~�9t 532t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 533t 61pw        sq ~��Z�pq ~ q ~�9t 533t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 534t 75pw        sq ~��Z�1q ~ q ~�9t 534t 84pw@M]��%��sq ~��Z�Pq ~ q ~�9t 535t 75pw        sq ~��Z��q ~ q ~�9t 535t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 536t 61pw        sq ~��Z��q ~ q ~�9t 536t 84pw@F�U�i�sq ~��Z�tq ~ q ~�9t 537t 84pw@F�U�i�sq ~��Z��q ~ q ~�9t 538t 75pw        sq ~��Z� 5q ~ q ~�9t 538t 84pw@5oz�G�sq ~��Z� Tq ~ q ~�9t 539t 75pw        sq ~��Z�#�q ~ q ~�9t 539t 84pw@5oz�G�sq ~��W�oq ~ q ~�9t 54t 18pw?����v�sq ~��W�J!q ~ q ~�9t 54t 5pw@4p$�Vn�sq ~��W�J@q ~ q ~�9t 54t 6pw        sq ~��Z�n�q ~ q ~�9t 540t 61pw        sq ~��Z�v�q ~ q ~�9t 540t 84pw@5oz�G�sq ~��Z�zMq ~ q ~�9t 541t 84pw@$      sq ~��Z�~q ~ q ~�9t 542t 84pw@5oz�G�sq ~��Z�y�q ~ q ~�9t 543t 61pw        sq ~��Z���q ~ q ~�9t 543t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 544t 75pw        sq ~��Z���q ~ q ~�9t 544t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 545t 75pw        sq ~��Z��Qq ~ q ~�9t 545t 84pw@5oz�G�sq ~��Z��3q ~ q ~�9t 546t 61pw        sq ~��Z��q ~ q ~�9t 546t 84pw@@�鹙�sq ~��Z��1q ~ q ~�9t 547t 75pw        sq ~��Z���q ~ q ~�9t 547t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 548t 61pw        sq ~��Z���q ~ q ~�9t 548t 84pw@$      sq ~��Z��Uq ~ q ~�9t 549t 84pw@F�U�i�sq ~��W�	�q ~ q ~�9t 55t 27pw@$      sq ~��Z���q ~ q ~�9t 550t 84pw@$      sq ~��Z��q ~ q ~�9t 551t 84pw@@�鹙�sq ~��Z��mq ~ q ~�9t 552t 84pw@$      sq ~��Z��q ~ q ~�9t 553t 75pw        sq ~��Z��.q ~ q ~�9t 553t 84pw@5oz�G�sq ~��Z��Mq ~ q ~�9t 554t 75pw        sq ~��Z���q ~ q ~�9t 554t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 555t 61pw        sq ~��Z���q ~ q ~�9t 555t 84pw@$      sq ~��Z�qq ~ q ~�9t 556t 84pw@$      sq ~��Z��q ~ q ~�9t 557t 75pw        sq ~��Z�2q ~ q ~�9t 557t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 558t 84pw@$      sq ~��Z��q ~ q ~�9t 559t 84pw@F�U�i�sq ~��W�6q ~ q ~�9t 56t 24pw@#�2�?sq ~��Z�[�q ~ q ~�9t 560t 75pw        sq ~��Z�_Jq ~ q ~�9t 560t 84pw@@�鹙�sq ~��Z�_iq ~ q ~�9t 561t 75pw        sq ~��Z�cq ~ q ~�9t 561t 84pw@$      sq ~��Z�f�q ~ q ~�9t 562t 84pw@@�鹙�sq ~��Z�f�q ~ q ~�9t 563t 75pw        sq ~��Z�j�q ~ q ~�9t 563t 84pw@5oz�G�sq ~��Z�foq ~ q ~�9t 564t 61pw        sq ~��Z�nNq ~ q ~�9t 564t 84pw@5oz�G�sq ~��Z�nmq ~ q ~�9t 565t 75pw        sq ~��Z�rq ~ q ~�9t 565t 84pw@5oz�G�sq ~��Z�r.q ~ q ~�9t 566t 75pw        sq ~��Z�u�q ~ q ~�9t 566t 84pw@5oz�G�sq ~��Z�y�q ~ q ~�9t 567t 84pw@@�鹙�sq ~��Z�y�q ~ q ~�9t 568t 75pw        sq ~��Z�}Rq ~ q ~�9t 568t 84pw@F�U�i�sq ~��Z�y4q ~ q ~�9t 569t 61pw        sq ~��Z��q ~ q ~�9t 569t 84pw@@�鹙�sq ~��W�q ~ q ~�9t 57t 13pw@$      sq ~��W�5q ~ q ~�9t 57t 26pw        sq ~��Z�өq ~ q ~�9t 570t 84pw@$      sq ~��Z���q ~ q ~�9t 571t 75pw        sq ~��Z��jq ~ q ~�9t 571t 84pw@5oz�G�sq ~��Z�׉q ~ q ~�9t 572t 75pw        sq ~��Z��+q ~ q ~�9t 572t 84pw@$      sq ~��Z��q ~ q ~�9t 573t 61pw        sq ~��Z���q ~ q ~�9t 573t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 574t 61pw        sq ~��Z��q ~ q ~�9t 574t 84pw@@�鹙�sq ~��Z��nq ~ q ~�9t 575t 84pw@@�鹙�sq ~��Z��/q ~ q ~�9t 576t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 577t 61pw        sq ~��Z���q ~ q ~�9t 577t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 578t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 579t 61pw        sq ~��Z��rq ~ q ~�9t 579t 84pw@$      sq ~��W�Tq ~ q ~�9t 58t 17pw@@w���Ӱsq ~��W��q ~ q ~�9t 58t 40pw@63�R���sq ~��W� wq ~ q ~�9t 58t 58pw        sq ~��Z�Hq ~ q ~�9t 580t 84pw@F�U�i�sq ~��Z�C�q ~ q ~�9t 581t 61pw        sq ~��Z�K�q ~ q ~�9t 581t 84pw@5oz�G�sq ~��Z�G�q ~ q ~�9t 582t 61pw        sq ~��Z�O�q ~ q ~�9t 582t 84pw@@�鹙�sq ~��Z�Klq ~ q ~�9t 583t 61pw        sq ~��Z�SKq ~ q ~�9t 583t 84pw@5oz�G�sq ~��Z�O-q ~ q ~�9t 584t 61pw        sq ~��Z�Wq ~ q ~�9t 584t 84pw@5oz�G�sq ~��Z�W+q ~ q ~�9t 585t 75pw        sq ~��Z�Z�q ~ q ~�9t 585t 84pw@5oz�G�sq ~��Z�Z�q ~ q ~�9t 586t 75pw        sq ~��Z�^�q ~ q ~�9t 586t 84pw@5oz�G�sq ~��Z�Zpq ~ q ~�9t 587t 61pw        sq ~��Z�bOq ~ q ~�9t 587t 84pw@$      sq ~��Z�bnq ~ q ~�9t 588t 75pw        sq ~��Z�fq ~ q ~�9t 588t 84pw@@�鹙�sq ~��Z�f/q ~ q ~�9t 589t 75pw        sq ~��Z�i�q ~ q ~�9t 589t 84pw@5oz�G�sq ~��W�yq ~ q ~�9t 59t 24pw�����sq ~��W��q ~ q ~�9t 59t 31pw@&j����sq ~��W�Yq ~ q ~�9t 59t 35pw        sq ~��Z���q ~ q ~�9t 590t 61pw        sq ~��Z��gq ~ q ~�9t 590t 84pw@F�U�i�sq ~��Z��Iq ~ q ~�9t 591t 61pw        sq ~��Z��(q ~ q ~�9t 591t 84pw@$      sq ~��Z��
q ~ q ~�9t 592t 61pw        sq ~��Z���q ~ q ~�9t 592t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 593t 61pw        sq ~��Z�Ǫq ~ q ~�9t 593t 84pw@5oz�G�sq ~��Z�Ìq ~ q ~�9t 594t 61pw        sq ~��Z��kq ~ q ~�9t 594t 84pw@@�鹙�sq ~��Z�ˊq ~ q ~�9t 595t 75pw        sq ~��Z��,q ~ q ~�9t 595t 84pw@$      sq ~��Z��Kq ~ q ~�9t 596t 75pw        sq ~��Z���q ~ q ~�9t 596t 84pw@$      sq ~��Z��q ~ q ~�9t 597t 75pw        sq ~��Z�֮q ~ q ~�9t 597t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 598t 75pw        sq ~��Z��oq ~ q ~�9t 598t 84pw@$      sq ~��Z�ڎq ~ q ~�9t 599t 75pw        sq ~��Z��0q ~ q ~�9t 599t 84pw@@�鹙�sq ~��W�9]q ~ q ~�9t 6t 0pw��!�8uLsq ~��W��Nq ~ q ~�9t 6t 10pw@#ӭRnx�sq ~��W��q ~ q ~�9t 6t 12pw�Ն��2sq ~��W��q ~ q ~�9t 6t 16pw@�J��rsq ~��W��Fq ~ q ~�9t 6t 18pw@.;PR�tsq ~��W��Mq ~ q ~�9t 6t 22pw��'Ek6Bsq ~��W��q ~ q ~�9t 6t 28pw?��RGD�sq ~��W��&q ~ q ~�9t 6t 29pw�uv���sq ~��W��q ~ q ~�9t 6t 32pw?��ҕ��usq ~��W���q ~ q ~�9t 6t 37pw��N�&sq ~��W��Kq ~ q ~�9t 6t 46pw?�PE"�sq ~��W�9�q ~ q ~�9t 6t 5pw?�C�ݓ�sq ~��W� qq ~ q ~�9t 6t 51pw@&p�<j#sq ~��W�:q ~ q ~�9t 6t 6pw@4�����vsq ~��W�gNq ~ q ~�9t 60t 14pw��+��k{sq ~��WƯ�q ~ q ~�9t 60t 8pw@$,[^��sq ~��Z���q ~ q ~�9t 600t 61pw        sq ~��Z���q ~ q ~�9t 600t 84pw@5oz�G�sq ~��Z��Rq ~ q ~�9t 601t 84pw@$      sq ~��Z��q ~ q ~�9t 602t 84pw@5oz�G�sq ~��Z��2q ~ q ~�9t 603t 75pw        sq ~��Z���q ~ q ~�9t 603t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 604t 75pw        sq ~��Z�˕q ~ q ~�9t 604t 84pw@5oz�G�sq ~��Z��Vq ~ q ~�9t 605t 84pw@5oz�G�sq ~��Z��8q ~ q ~�9t 606t 61pw        sq ~��Z��q ~ q ~�9t 606t 84pw@@�鹙�sq ~��Z��6q ~ q ~�9t 607t 75pw        sq ~��Z���q ~ q ~�9t 607t 84pw@$      sq ~��Z�Һq ~ q ~�9t 608t 61pw        sq ~��Z�ڙq ~ q ~�9t 608t 84pw@@�鹙�sq ~��Z��Zq ~ q ~�9t 609t 84pw@@�鹙�sq ~��W�kq ~ q ~�9t 61t 14pw@ i��|�Rsq ~��W�k.q ~ q ~�9t 61t 15pw@�mᔫ�sq ~��W�nTq ~ q ~�9t 61t 20pw        sq ~��WƳ�q ~ q ~�9t 61t 9pw?���}!x�sq ~��Z�0�q ~ q ~�9t 610t 84pw@5oz�G�sq ~��Z�,�q ~ q ~�9t 611t 61pw        sq ~��Z�4�q ~ q ~�9t 611t 84pw@F�U�i�sq ~��Z�0�q ~ q ~�9t 612t 61pw        sq ~��Z�8rq ~ q ~�9t 612t 84pw@5oz�G�sq ~��Z�<3q ~ q ~�9t 613t 84pw@$      sq ~��Z�<Rq ~ q ~�9t 614t 75pw        sq ~��Z�?�q ~ q ~�9t 614t 84pw@$      sq ~��Z�;�q ~ q ~�9t 615t 61pw        sq ~��Z�C�q ~ q ~�9t 615t 84pw@$      sq ~��Z�Gvq ~ q ~�9t 616t 84pw@$      sq ~��Z�K7q ~ q ~�9t 617t 84pw@$      sq ~��Z�N�q ~ q ~�9t 618t 84pw@@�鹙�sq ~��Z�Oq ~ q ~�9t 619t 75pw        sq ~��Z�R�q ~ q ~�9t 619t 84pw@@�鹙�sq ~��W�n�q ~ q ~�9t 62t 14pw@L��X~sq ~��W�n�q ~ q ~�9t 62t 15pw��"��۹sq ~��W�rq ~ q ~�9t 62t 20pw        sq ~��Wǅq ~ q ~�9t 62t 72pw���� 1�sq ~��WƷ[q ~ q ~�9t 62t 8pw@\<�HNsq ~��WƷzq ~ q ~�9t 62t 9pw��7D��dsq ~��Z��Oq ~ q ~�9t 620t 84pw@F�U�i�sq ~��Z��1q ~ q ~�9t 621t 61pw        sq ~��Z��q ~ q ~�9t 621t 84pw@$      sq ~��Z���q ~ q ~�9t 622t 61pw        sq ~��Z���q ~ q ~�9t 622t 84pw@$      sq ~��Z���q ~ q ~�9t 623t 61pw        sq ~��Z���q ~ q ~�9t 623t 84pw@5oz�G�sq ~��Z��Sq ~ q ~�9t 624t 84pw@5oz�G�sq ~��Z��rq ~ q ~�9t 625t 75pw        sq ~��Z��q ~ q ~�9t 625t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 626t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 627t 61pw        sq ~��Z���q ~ q ~�9t 627t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 628t 75pw        sq ~��Z��Wq ~ q ~�9t 628t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 629t 84pw@@�鹙�sq ~��WƺCq ~ q ~�9t 63t 1pw@&�'w�sq ~��Wǅq ~ q ~�9t 63t 62pw        sq ~��Z�q ~ q ~�9t 630t 75pw        sq ~��Z��q ~ q ~�9t 630t 84pw@@�鹙�sq ~��Z�oq ~ q ~�9t 631t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 632t 75pw        sq ~��Z�!0q ~ q ~�9t 632t 84pw@@�鹙�sq ~��Z�!Oq ~ q ~�9t 633t 75pw        sq ~��Z�$�q ~ q ~�9t 633t 84pw@5oz�G�sq ~��Z� �q ~ q ~�9t 634t 61pw        sq ~��Z�(�q ~ q ~�9t 634t 84pw@5oz�G�sq ~��Z�(�q ~ q ~�9t 635t 75pw        sq ~��Z�,sq ~ q ~�9t 635t 84pw@F�U�i�sq ~��Z�(Uq ~ q ~�9t 636t 61pw        sq ~��Z�04q ~ q ~�9t 636t 84pw@$      sq ~��Z�,q ~ q ~�9t 637t 61pw        sq ~��Z�3�q ~ q ~�9t 637t 84pw@@�鹙�sq ~��Z�7�q ~ q ~�9t 638t 84pw@@�鹙�sq ~��Z�7�q ~ q ~�9t 639t 75pw        sq ~��Z�;wq ~ q ~�9t 639t 84pw@$      sq ~��W�~q ~ q ~�9t 64t 36pw        sq ~��Wƾaq ~ q ~�9t 64t 4pw@5oz�G�sq ~��Wǅ�q ~ q ~�9t 64t 59pw@5oz�G�sq ~��Z��.q ~ q ~�9t 640t 61pw        sq ~��Z��q ~ q ~�9t 640t 84pw@$      sq ~��Z���q ~ q ~�9t 641t 61pw        sq ~��Z���q ~ q ~�9t 641t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 642t 61pw        sq ~��Z���q ~ q ~�9t 642t 84pw@$      sq ~��Z��Pq ~ q ~�9t 643t 84pw@5oz�G�sq ~��Z��2q ~ q ~�9t 644t 61pw        sq ~��Z��q ~ q ~�9t 644t 84pw@5oz�G�sq ~��Z��0q ~ q ~�9t 645t 75pw        sq ~��Z���q ~ q ~�9t 645t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 646t 75pw        sq ~��Z���q ~ q ~�9t 646t 84pw@5oz�G�sq ~��Z��uq ~ q ~�9t 647t 61pw        sq ~��Z��Tq ~ q ~�9t 647t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 648t 84pw@5oz�G�sq ~��Z��4q ~ q ~�9t 649t 75pw        sq ~��Z���q ~ q ~�9t 649t 84pw@5oz�G�sq ~��W�y�q ~ q ~�9t 65t 13pw        sq ~��W�}wq ~ q ~�9t 65t 21pw@/j�ysq ~��W��"q ~ q ~�9t 65t 4pw�p��N1 �sq ~��WǅVq ~ q ~�9t 65t 44pw���-k��sq ~��Wǅuq ~ q ~�9t 65t 45pw@1���ϑ�sq ~��Wǉ�q ~ q ~�9t 65t 59pw�3��m��sq ~��Z�lq ~ q ~�9t 650t 84pw@5oz�G�sq ~��Z��Nq ~ q ~�9t 651t 61pw        sq ~��Z�-q ~ q ~�9t 651t 84pw@5oz�G�sq ~��Z�	�q ~ q ~�9t 652t 84pw@5oz�G�sq ~��Z�
q ~ q ~�9t 653t 75pw        sq ~��Z��q ~ q ~�9t 653t 84pw@$      sq ~��Z�pq ~ q ~�9t 654t 84pw@5oz�G�sq ~��Z�1q ~ q ~�9t 655t 84pw@5oz�G�sq ~��Z�Pq ~ q ~�9t 656t 75pw        sq ~��Z��q ~ q ~�9t 656t 84pw@@�鹙�sq ~��Z�q ~ q ~�9t 657t 75pw        sq ~��Z��q ~ q ~�9t 657t 84pw@$      sq ~��Z��q ~ q ~�9t 658t 61pw        sq ~��Z� tq ~ q ~�9t 658t 84pw@@�鹙�sq ~��Z�$5q ~ q ~�9t 659t 84pw@@�鹙�sq ~��Wǁ�q ~ q ~�9t 66t 25pw        sq ~��WǍTq ~ q ~�9t 66t 58pw@5oz�G�sq ~��WǑ4q ~ q ~�9t 66t 69pw@5oz�G�sq ~��WǓ�q ~ q ~�9t 66t 70pw        sq ~��Z�s)q ~ q ~�9t 660t 75pw        sq ~��Z�v�q ~ q ~�9t 660t 84pw@@�鹙�sq ~��Z�r�q ~ q ~�9t 661t 61pw        sq ~��Z�z�q ~ q ~�9t 661t 84pw@5oz�G�sq ~��Z�~Mq ~ q ~�9t 662t 84pw@$      sq ~��Z��q ~ q ~�9t 663t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 664t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 665t 61pw        sq ~��Z���q ~ q ~�9t 665t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 666t 75pw        sq ~��Z��Qq ~ q ~�9t 666t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 667t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 668t 61pw        sq ~��Z���q ~ q ~�9t 668t 84pw@$      sq ~��Z���q ~ q ~�9t 669t 84pw@$      sq ~��WǄ�q ~ q ~�9t 67t 21pw@!�_��sq ~��Wǌ�q ~ q ~�9t 67t 44pw@�g��sq ~��Wǌ�q ~ q ~�9t 67t 45pw@$�ܮ��sq ~��WǑ4q ~ q ~�9t 67t 59pw��i���sq ~��Z��q ~ q ~�9t 670t 75pw        sq ~��Z��*q ~ q ~�9t 670t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 671t 61pw        sq ~��Z���q ~ q ~�9t 671t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 672t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 673t 61pw        sq ~��Z��mq ~ q ~�9t 673t 84pw@@�鹙�sq ~��Z��Oq ~ q ~�9t 674t 61pw        sq ~��Z��.q ~ q ~�9t 674t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 675t 61pw        sq ~��Z���q ~ q ~�9t 675t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 676t 61pw        sq ~��Z��q ~ q ~�9t 676t 84pw@5oz�G�sq ~��Z�qq ~ q ~�9t 677t 84pw@5oz�G�sq ~��Z�Sq ~ q ~�9t 678t 61pw        sq ~��Z�	2q ~ q ~�9t 678t 84pw@5oz�G�sq ~��Z�q ~ q ~�9t 679t 61pw        sq ~��Z��q ~ q ~�9t 679t 84pw@@�鹙�sq ~��WǅVq ~ q ~�9t 68t 14pw@!�d_/�sq ~��Wǅuq ~ q ~�9t 68t 15pw�h��Wsq ~��Wǐzq ~ q ~�9t 68t 43pw�����sq ~��WǛ�q ~ q ~�9t 68t 72pw        sq ~��W���q ~ q ~�9t 68t 8pw@+�6�t��sq ~��Z�[�q ~ q ~�9t 680t 75pw        sq ~��Z�_�q ~ q ~�9t 680t 84pw@$      sq ~��Z�cJq ~ q ~�9t 681t 84pw@$      sq ~��Z�gq ~ q ~�9t 682t 84pw@@�鹙�sq ~��Z�j�q ~ q ~�9t 683t 84pw@$      sq ~��Z�n�q ~ q ~�9t 684t 84pw@@�鹙�sq ~��Z�rNq ~ q ~�9t 685t 84pw@@�鹙�sq ~��Z�rmq ~ q ~�9t 686t 75pw        sq ~��Z�vq ~ q ~�9t 686t 84pw@5oz�G�sq ~��Z�q�q ~ q ~�9t 687t 61pw��3��sq ~��Z�y�q ~ q ~�9t 687t 84pw@6fΪ/|ksq ~��Z�}�q ~ q ~�9t 688t 84pw@@�鹙�sq ~��Z��Rq ~ q ~�9t 689t 84pw@5oz�G�sq ~��Wǌ�q ~ q ~�9t 69t 24pw�+��E٧sq ~��Wǐ<q ~ q ~�9t 69t 31pw@'���	�Gsq ~��Wǜ9q ~ q ~�9t 69t 67pw        sq ~��Wǟ�q ~ q ~�9t 69t 76pw@$      sq ~��Z���q ~ q ~�9t 690t 84pw@$      sq ~��Z���q ~ q ~�9t 691t 61pw        sq ~��Z�שq ~ q ~�9t 691t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 692t 75pw        sq ~��Z��jq ~ q ~�9t 692t 84pw@5oz�G�sq ~��Z��+q ~ q ~�9t 693t 84pw@$      sq ~��Z���q ~ q ~�9t 694t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 695t 75pw        sq ~��Z��q ~ q ~�9t 695t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 696t 61pw        sq ~��Z��nq ~ q ~�9t 696t 84pw@5oz�G�sq ~��Z��/q ~ q ~�9t 697t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 698t 61pw        sq ~��Z���q ~ q ~�9t 698t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 699t 75pw        sq ~��Z���q ~ q ~�9t 699t 84pw@$      sq ~��W� qq ~ q ~�9t 7t 41pw@'�.��R�sq ~��W�>q ~ q ~�9t 7t 8pw        sq ~��W�>5q ~ q ~�9t 7t 9pw        sq ~��W���q ~ q ~�9t 70t 55pw@@�鹙�sq ~��Z��q ~ q ~�9t 700t 84pw@F�U�i�sq ~��Z��1q ~ q ~�9t 701t 75pw        sq ~��Z���q ~ q ~�9t 701t 84pw@$      sq ~��Z�۔q ~ q ~�9t 702t 84pw@5oz�G�sq ~��Z�۳q ~ q ~�9t 703t 75pw        sq ~��Z��Uq ~ q ~�9t 703t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 704t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 705t 61pw        sq ~��Z���q ~ q ~�9t 705t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 706t 75pw        sq ~��Z��q ~ q ~�9t 706t 84pw@$      sq ~��Z��zq ~ q ~�9t 707t 61pw        sq ~��Z��Yq ~ q ~�9t 707t 84pw@@�鹙�sq ~��Z��;q ~ q ~�9t 708t 61pw        sq ~��Z��q ~ q ~�9t 708t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 709t 61pw        sq ~��Z���q ~ q ~�9t 709t 84pw@@�鹙�sq ~��W��q ~ q ~�9t 71t 43pw        sq ~��W���q ~ q ~�9t 71t 72pw@$      sq ~��Z�@�q ~ q ~�9t 710t 61pw        sq ~��Z�Hqq ~ q ~�9t 710t 84pw@5oz�G�sq ~��Z�L2q ~ q ~�9t 711t 84pw@@�鹙�sq ~��Z�O�q ~ q ~�9t 712t 84pw@$      sq ~��Z�K�q ~ q ~�9t 713t 61pw        sq ~��Z�S�q ~ q ~�9t 713t 84pw@5oz�G�sq ~��Z�Wuq ~ q ~�9t 714t 84pw@5oz�G�sq ~��Z�SWq ~ q ~�9t 715t 61pw        sq ~��Z�[6q ~ q ~�9t 715t 84pw@$      sq ~��Z�^�q ~ q ~�9t 716t 84pw@F�U�i�sq ~��Z�Z�q ~ q ~�9t 717t 61pw        sq ~��Z�b�q ~ q ~�9t 717t 84pw@5oz�G�sq ~��Z�fyq ~ q ~�9t 718t 84pw@$      sq ~��Z�f�q ~ q ~�9t 719t 75pw        sq ~��Z�j:q ~ q ~�9t 719t 84pw@5oz�G�sq ~��W��Rq ~ q ~�9t 72t 55pw        sq ~��W���q ~ q ~�9t 72t 73pw@$      sq ~��Z̹.q ~ q ~�9t 720t 75pw        sq ~��Z̼�q ~ q ~�9t 720t 84pw@5oz�G�sq ~��Z̼�q ~ q ~�9t 721t 75pw        sq ~��Z���q ~ q ~�9t 721t 84pw@F�U�i�sq ~��Z��Rq ~ q ~�9t 722t 84pw@F�U�i�sq ~��Z��4q ~ q ~�9t 723t 61pw        sq ~��Z��q ~ q ~�9t 723t 84pw@$      sq ~��Z��2q ~ q ~�9t 724t 75pw        sq ~��Z���q ~ q ~�9t 724t 84pw@5oz�G�sq ~��Z�Ƕq ~ q ~�9t 725t 61pw        sq ~��Z�ϕq ~ q ~�9t 725t 84pw@@�鹙�sq ~��Z��wq ~ q ~�9t 726t 61pw        sq ~��Z��Vq ~ q ~�9t 726t 84pw@@�鹙�sq ~��Z��uq ~ q ~�9t 727t 75pw        sq ~��Z��q ~ q ~�9t 727t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 728t 61pw        sq ~��Z���q ~ q ~�9t 728t 84pw@$      sq ~��Z�ֺq ~ q ~�9t 729t 61pw        sq ~��Z�ޙq ~ q ~�9t 729t 84pw@@�鹙�sq ~��W��2q ~ q ~�9t 73t 56pw@$      sq ~��W��vq ~ q ~�9t 73t 74pw@$      sq ~��Z�1/q ~ q ~�9t 730t 84pw@$      sq ~��Z�4�q ~ q ~�9t 731t 84pw@@�鹙�sq ~��Z�8�q ~ q ~�9t 732t 84pw@5oz�G�sq ~��Z�4�q ~ q ~�9t 733t 61pw        sq ~��Z�<rq ~ q ~�9t 733t 84pw@@�鹙�sq ~��Z�<�q ~ q ~�9t 734t 75pw        sq ~��Z�@3q ~ q ~�9t 734t 84pw@$      sq ~��Z�@Rq ~ q ~�9t 735t 75pw        sq ~��Z�C�q ~ q ~�9t 735t 84pw@5oz�G�sq ~��Z�?�q ~ q ~�9t 736t 61pw        sq ~��Z�G�q ~ q ~�9t 736t 84pw@#��Ё�sq ~��Z�Kvq ~ q ~�9t 737t 84pw@F�U�i�sq ~��Z�O7q ~ q ~�9t 738t 84pw@$      sq ~��Z�R�q ~ q ~�9t 739t 84pw@#ٳ�:�sq ~��W��q ~ q ~�9t 74t 14pw����|�ɵsq ~��W���q ~ q ~�9t 74t 15pw@U}�D��sq ~��W���q ~ q ~�9t 74t 43pw        sq ~��W� �q ~ q ~�9t 74t 72pw�����P�sq ~��W�3[q ~ q ~�9t 74t 9pw?���	9�~sq ~��Z͝�q ~ q ~�9t 740t 61pw        sq ~��Zͥ�q ~ q ~�9t 740t 84pw@@�鹙�sq ~��Zͥ�q ~ q ~�9t 741t 75pw        sq ~��ZͩOq ~ q ~�9t 741t 84pw@$      sq ~��Zͥ1q ~ q ~�9t 742t 61pw        sq ~��Zͭq ~ q ~�9t 742t 84pw@@�鹙�sq ~��Zͨ�q ~ q ~�9t 743t 61pw        sq ~��ZͰ�q ~ q ~�9t 743t 84pw@$      sq ~��Zʹ�q ~ q ~�9t 744t 84pw@@�鹙�sq ~��Zʹ�q ~ q ~�9t 745t 75pw        sq ~��Z͸Sq ~ q ~�9t 745t 84pw@@�鹙�sq ~��Zʹ5q ~ q ~�9t 746t 61pw        sq ~��Zͼq ~ q ~�9t 746t 84pw@@�鹙�sq ~��ZͿ�q ~ q ~�9t 747t 84pw@5oz�G�sq ~��ZͿ�q ~ q ~�9t 748t 75pw        sq ~��Z�Öq ~ q ~�9t 748t 84pw@$      sq ~��Z�õq ~ q ~�9t 749t 75pw        sq ~��Z��Wq ~ q ~�9t 749t 84pw@5oz�G�sq ~��W��q ~ q ~�9t 75t 27pw@)ꑷ(�lsq ~��W� �q ~ q ~�9t 75t 60pw        sq ~��Z�q ~ q ~�9t 750t 61pw        sq ~��Z��q ~ q ~�9t 750t 84pw@$      sq ~��Z��q ~ q ~�9t 751t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 752t 75pw        sq ~��Z�!oq ~ q ~�9t 752t 84pw@5oz�G�sq ~��Z�!�q ~ q ~�9t 753t 75pw        sq ~��Z�%0q ~ q ~�9t 753t 84pw@5oz�G�sq ~��Z�(�q ~ q ~�9t 754t 84pw@$      sq ~��Z�,�q ~ q ~�9t 755t 84pw@$      sq ~��Z�0sq ~ q ~�9t 756t 84pw@$      sq ~��Z�,Uq ~ q ~�9t 757t 61pw        sq ~��Z�44q ~ q ~�9t 757t 84pw@$      sq ~��Z�4Sq ~ q ~�9t 758t 75pw        sq ~��Z�7�q ~ q ~�9t 758t 84pw@@�鹙�sq ~��Z�8q ~ q ~�9t 759t 75pw        sq ~��Z�;�q ~ q ~�9t 759t 84pw@5oz�G�sq ~��W��q ~ q ~�9t 76t 61pw        sq ~��W��q ~ q ~�9t 76t 75pw@@�鹙�sq ~��ZΎLq ~ q ~�9t 760t 84pw@5oz�G�sq ~��ZΊ.q ~ q ~�9t 761t 61pw        sq ~��ZΒq ~ q ~�9t 761t 84pw@$      sq ~��Z΍�q ~ q ~�9t 762t 61pw        sq ~��ZΕ�q ~ q ~�9t 762t 84pw@$      sq ~��ZΑ�q ~ q ~�9t 763t 61pw        sq ~��ZΙ�q ~ q ~�9t 763t 84pw@5oz�G�sq ~��ZΕqq ~ q ~�9t 764t 61pw        sq ~��ZΝPq ~ q ~�9t 764t 84pw@$      sq ~��ZΡq ~ q ~�9t 765t 84pw@$      sq ~��ZΤ�q ~ q ~�9t 766t 84pw@5oz�G�sq ~��ZΨ�q ~ q ~�9t 767t 84pw@$      sq ~��ZΨ�q ~ q ~�9t 768t 75pw        sq ~��ZάTq ~ q ~�9t 768t 84pw@F�U�i�sq ~��Zάsq ~ q ~�9t 769t 75pw        sq ~��Zΰq ~ q ~�9t 769t 84pw@5oz�G�sq ~��W���q ~ q ~�9t 77t 14pw��x�,���sq ~��W��q ~ q ~�9t 77t 15pw���"A�sq ~��W�>q ~ q ~�9t 77t 8pw        sq ~��W�>�q ~ q ~�9t 77t 9pw@#>=���sq ~��Z��q ~ q ~�9t 770t 84pw@@�鹙�sq ~��Z�lq ~ q ~�9t 771t 84pw@5oz�G�sq ~��Z�Nq ~ q ~�9t 772t 61pw        sq ~��Z�
-q ~ q ~�9t 772t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 773t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 774t 84pw@$      sq ~��Z�pq ~ q ~�9t 775t 84pw@@�鹙�sq ~��Z�1q ~ q ~�9t 776t 84pw@5oz�G�sq ~��Z�Pq ~ q ~�9t 777t 75pw        sq ~��Z��q ~ q ~�9t 777t 84pw@@�鹙�sq ~��Z� �q ~ q ~�9t 778t 84pw@F�U�i�sq ~��Z��q ~ q ~�9t 779t 61pw        sq ~��Z�$tq ~ q ~�9t 779t 84pw@5oz�G�sq ~��W��q ~ q ~�9t 78t 56pw@$      sq ~��W�;q ~ q ~�9t 78t 74pw@$      sq ~��Z�shq ~ q ~�9t 780t 75pw        sq ~��Z�w
q ~ q ~�9t 780t 84pw@F�U�i�sq ~��Z�z�q ~ q ~�9t 781t 84pw@@�鹙�sq ~��Z�z�q ~ q ~�9t 782t 75pw        sq ~��Z�~�q ~ q ~�9t 782t 84pw@5oz�G�sq ~��Z�znq ~ q ~�9t 783t 61pw        sq ~��ZςMq ~ q ~�9t 783t 84pw@$      sq ~��Zςlq ~ q ~�9t 784t 75pw        sq ~��Zφq ~ q ~�9t 784t 84pw@@�鹙�sq ~��Zφ-q ~ q ~�9t 785t 75pw        sq ~��Zω�q ~ q ~�9t 785t 84pw@5oz�G�sq ~��Zύ�q ~ q ~�9t 786t 84pw@5oz�G�sq ~��Zωrq ~ q ~�9t 787t 61pw        sq ~��ZϑQq ~ q ~�9t 787t 84pw@@�鹙�sq ~��Zϑpq ~ q ~�9t 788t 75pw        sq ~��Zϕq ~ q ~�9t 788t 84pw@F�U�i�sq ~��ZϘ�q ~ q ~�9t 789t 84pw@5oz�G�sq ~��W�E(q ~ q ~�9t 79t 1pw@#�^e�R�sq ~��W��q ~ q ~�9t 79t 62pw@$      sq ~��Z��q ~ q ~�9t 790t 61pw        sq ~��Z��iq ~ q ~�9t 790t 84pw@5oz�G�sq ~��Z��*q ~ q ~�9t 791t 84pw@$      sq ~��Z��Iq ~ q ~�9t 792t 75pw        sq ~��Z���q ~ q ~�9t 792t 84pw@$      sq ~��Z���q ~ q ~�9t 793t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 794t 61pw        sq ~��Z��mq ~ q ~�9t 794t 84pw@$      sq ~��Z��.q ~ q ~�9t 795t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 796t 61pw        sq ~��Z��q ~ q ~�9t 796t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 797t 61pw        sq ~��Z��q ~ q ~�9t 797t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 798t 75pw        sq ~��Z�	qq ~ q ~�9t 798t 84pw@5oz�G�sq ~��Z�	�q ~ q ~�9t 799t 75pw        sq ~��Z�2q ~ q ~�9t 799t 84pw@$      sq ~��W���q ~ q ~�9t 8t 10pw        sq ~��W��q ~ q ~�9t 8t 46pw@5oz�G�sq ~��W�b�q ~ q ~�9t 80t 64pw@5oz�G�sq ~��Z���q ~ q ~�9t 800t 75pw        sq ~��Z��q ~ q ~�9t 800t 84pw@$      sq ~��Z��uq ~ q ~�9t 801t 61pw        sq ~��Z��Tq ~ q ~�9t 801t 84pw@$      sq ~��Z��sq ~ q ~�9t 802t 75pw        sq ~��Z��q ~ q ~�9t 802t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 803t 61pw        sq ~��Z���q ~ q ~�9t 803t 84pw@$>�(R=�sq ~��Z���q ~ q ~�9t 804t 75pw        sq ~��Z���q ~ q ~�9t 804t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 805t 75pw        sq ~��Z��Xq ~ q ~�9t 805t 84pw@5oz�G�sq ~��Z��:q ~ q ~�9t 806t 61pw        sq ~��Z�q ~ q ~�9t 806t 84pw@F�U�i�sq ~��Z��q ~ q ~�9t 807t 84pw@$      sq ~��Z�	�q ~ q ~�9t 808t 84pw@$      sq ~��Z�}q ~ q ~�9t 809t 61pw        sq ~��Z�\q ~ q ~�9t 809t 84pw@@�鹙�sq ~��W�[0q ~ q ~�9t 81t 33pw@$      sq ~��W�f�q ~ q ~�9t 81t 65pw        sq ~��Z�\Pq ~ q ~�9t 810t 75pw        sq ~��Z�_�q ~ q ~�9t 810t 84pw@@�鹙�sq ~��Z�`q ~ q ~�9t 811t 75pw        sq ~��Z�c�q ~ q ~�9t 811t 84pw@@�鹙�sq ~��Z�c�q ~ q ~�9t 812t 75pw        sq ~��Z�gtq ~ q ~�9t 812t 84pw@$      sq ~��Z�k5q ~ q ~�9t 813t 84pw@@�鹙�sq ~��Z�n�q ~ q ~�9t 814t 84pw@$      sq ~��Z�j�q ~ q ~�9t 815t 61pw        sq ~��Z�r�q ~ q ~�9t 815t 84pw@5���Q�sq ~��Z�vxq ~ q ~�9t 816t 84pw@$      sq ~��Z�v�q ~ q ~�9t 817t 75pw        sq ~��Z�z9q ~ q ~�9t 817t 84pw@@�鹙�sq ~��Z�zXq ~ q ~�9t 818t 75pw        sq ~��Z�}�q ~ q ~�9t 818t 84pw@5oz�G�sq ~��Z�~q ~ q ~�9t 819t 75pw        sq ~��Zځ�q ~ q ~�9t 819t 84pw@$      sq ~��W�[nq ~ q ~�9t 82t 25pw        sq ~��W�gq ~ q ~�9t 82t 58pw@$      sq ~��W�j�q ~ q ~�9t 82t 69pw@$      sq ~��Z�Яq ~ q ~�9t 820t 75pw        sq ~��Z��Qq ~ q ~�9t 820t 84pw@5oz�G�sq ~��Z��pq ~ q ~�9t 821t 75pw        sq ~��Z��q ~ q ~�9t 821t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 822t 61pw        sq ~��Z���q ~ q ~�9t 822t 84pw@@�鹙�sq ~��Z�ߔq ~ q ~�9t 823t 84pw@5oz�G�sq ~��Z��Uq ~ q ~�9t 824t 84pw@5oz�G�sq ~��Z��tq ~ q ~�9t 825t 75pw        sq ~��Z��q ~ q ~�9t 825t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 826t 61pw        sq ~��Z���q ~ q ~�9t 826t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 827t 75pw        sq ~��Z��q ~ q ~�9t 827t 84pw@$      sq ~��Z��zq ~ q ~�9t 828t 61pw        sq ~��Z��Yq ~ q ~�9t 828t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 829t 84pw@5oz�G�sq ~��W�_/q ~ q ~�9t 83t 25pw�F�~V��sq ~��W�bUq ~ q ~�9t 83t 30pw@%��/�Hsq ~��W�j�q ~ q ~�9t 83t 57pw@%���(�sq ~��Z�@�q ~ q ~�9t 830t 61pw        sq ~��Z�H�q ~ q ~�9t 830t 84pw@6��Dڠsq ~��Z�H�q ~ q ~�9t 831t 75pw        sq ~��Z�Lqq ~ q ~�9t 831t 84pw@5oz�G�sq ~��Z�P2q ~ q ~�9t 832t 84pw@5oz�G�sq ~��Z�PQq ~ q ~�9t 833t 75pw        sq ~��Z�S�q ~ q ~�9t 833t 84pw@F�U�i�sq ~��Z�W�q ~ q ~�9t 834t 84pw@5oz�G�sq ~��Z�[uq ~ q ~�9t 835t 84pw@$      sq ~��Z�_6q ~ q ~�9t 836t 84pw@$      sq ~��Z�[q ~ q ~�9t 837t 61pw        sq ~��Z�b�q ~ q ~�9t 837t 84pw@5oz�G�sq ~��Z�cq ~ q ~�9t 838t 75pw        sq ~��Z�f�q ~ q ~�9t 838t 84pw@@�鹙�sq ~��Z�f�q ~ q ~�9t 839t 75pw        sq ~��Z�jyq ~ q ~�9t 839t 84pw@@�鹙�sq ~��WǦ�q ~ q ~�9t 84t 1pw@$e{i�sq ~��W�rq ~ q ~�9t 84t 66pw        sq ~��Z۵0q ~ q ~�9t 840t 61pw        sq ~��Z۽q ~ q ~�9t 840t 84pw@$      sq ~��Z���q ~ q ~�9t 841t 84pw@$      sq ~��Zۼ�q ~ q ~�9t 842t 61pw        sq ~��Z�đq ~ q ~�9t 842t 84pw@5oz�G�sq ~��Z�İq ~ q ~�9t 843t 75pw        sq ~��Z��Rq ~ q ~�9t 843t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 844t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 845t 61pw        sq ~��Z���q ~ q ~�9t 845t 84pw@F�U�i�sq ~��Z���q ~ q ~�9t 846t 75pw        sq ~��Z�ӕq ~ q ~�9t 846t 84pw@$      sq ~��Z��wq ~ q ~�9t 847t 61pw        sq ~��Z��Vq ~ q ~�9t 847t 84pw@5oz�G�sq ~��Z��uq ~ q ~�9t 848t 75pw        sq ~��Z��q ~ q ~�9t 848t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 849t 61pw        sq ~��Z���q ~ q ~�9t 849t 84pw@5oz�G�sq ~��W�rq ~ q ~�9t 85t 56pw@5oz�G�sq ~��W�yWq ~ q ~�9t 85t 74pw@5oz�G�sq ~��Z�-�q ~ q ~�9t 850t 75pw        sq ~��Z�1nq ~ q ~�9t 850t 84pw@$      sq ~��Z�5/q ~ q ~�9t 851t 84pw@"��r
sq ~��Z�5Nq ~ q ~�9t 852t 75pw        sq ~��Z�8�q ~ q ~�9t 852t 84pw@$      sq ~��Z�4�q ~ q ~�9t 853t 61pw        sq ~��Z�<�q ~ q ~�9t 853t 84pw@@�鹙�sq ~��Z�8�q ~ q ~�9t 854t 61pw        sq ~��Z�@rq ~ q ~�9t 854t 84pw@$      sq ~��Z�<Tq ~ q ~�9t 855t 61pw        sq ~��Z�D3q ~ q ~�9t 855t 84pw@5oz�G�sq ~��Z�G�q ~ q ~�9t 856t 84pw@"��a�5sq ~��Z�C�q ~ q ~�9t 857t 61pw        sq ~��Z�K�q ~ q ~�9t 857t 84pw@5oz�G�sq ~��Z�K�q ~ q ~�9t 858t 75pw        sq ~��Z�Ovq ~ q ~�9t 858t 84pw@5oz�G�sq ~��Z�O�q ~ q ~�9t 859t 75pw        sq ~��Z�S7q ~ q ~�9t 859t 84pw@@�鹙�sq ~��W�j�q ~ q ~�9t 86t 27pw@2ڐ��?sq ~��W�y�q ~ q ~�9t 86t 68pw        sq ~��Zܥ�q ~ q ~�9t 860t 84pw@@�鹙�sq ~��Zܡ�q ~ q ~�9t 861t 61pw        sq ~��Zܩ�q ~ q ~�9t 861t 84pw@5oz�G�sq ~��Zܥpq ~ q ~�9t 862t 61pw        sq ~��ZܭOq ~ q ~�9t 862t 84pw@$      sq ~��Zܩ1q ~ q ~�9t 863t 61pw        sq ~��Zܱq ~ q ~�9t 863t 84pw@#�B5_Z�sq ~��Zܴ�q ~ q ~�9t 864t 84pw@@�鹙�sq ~��Zܴ�q ~ q ~�9t 865t 75pw        sq ~��Zܸ�q ~ q ~�9t 865t 84pw@$      sq ~��ZܼSq ~ q ~�9t 866t 84pw@@�鹙�sq ~��Zܼrq ~ q ~�9t 867t 75pw        sq ~��Z��q ~ q ~�9t 867t 84pw@5oz�G�sq ~��Zܻ�q ~ q ~�9t 868t 61pw        sq ~��Z���q ~ q ~�9t 868t 84pw@$      sq ~��Zܿ�q ~ q ~�9t 869t 61pw        sq ~��Z�ǖq ~ q ~�9t 869t 84pw@F�U�i�sq ~��W�y8q ~ q ~�9t 87t 53pw        sq ~��W�yWq ~ q ~�9t 87t 54pw@5oz�G�sq ~��Z�Mq ~ q ~�9t 870t 61pw        sq ~��Z�,q ~ q ~�9t 870t 84pw@@�鹙�sq ~��Z�Kq ~ q ~�9t 871t 75pw        sq ~��Z��q ~ q ~�9t 871t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 872t 61pw        sq ~��Z�!�q ~ q ~�9t 872t 84pw@5oz�G�sq ~��Z�%oq ~ q ~�9t 873t 84pw@@�鹙�sq ~��Z�!Qq ~ q ~�9t 874t 61pw        sq ~��Z�)0q ~ q ~�9t 874t 84pw@@�鹙�sq ~��Z�,�q ~ q ~�9t 875t 84pw@5oz�G�sq ~��Z�-q ~ q ~�9t 876t 75pw        sq ~��Z�0�q ~ q ~�9t 876t 84pw@5oz�G�sq ~��Z�0�q ~ q ~�9t 877t 75pw        sq ~��Z�4sq ~ q ~�9t 877t 84pw@5oz�G�sq ~��Z�4�q ~ q ~�9t 878t 75pw        sq ~��Z�84q ~ q ~�9t 878t 84pw@5oz�G�sq ~��Z�8Sq ~ q ~�9t 879t 75pw        sq ~��Z�;�q ~ q ~�9t 879t 84pw@F�U�i�sq ~��W�nq ~ q ~�9t 88t 14pw@(0�!�sq ~��W�n3q ~ q ~�9t 88t 15pw���ۃ��sq ~��W�x�q ~ q ~�9t 88t 41pw���q{�sq ~��W�y8q ~ q ~�9t 88t 43pw        sq ~��Z݆�q ~ q ~�9t 880t 61pw        sq ~��Zݎ�q ~ q ~�9t 880t 84pw@@�鹙�sq ~��Zݎ�q ~ q ~�9t 881t 75pw        sq ~��ZݒLq ~ q ~�9t 881t 84pw@@�鹙�sq ~��Zݒkq ~ q ~�9t 882t 75pw        sq ~��Zݖq ~ q ~�9t 882t 84pw@$      sq ~��Zݙ�q ~ q ~�9t 883t 84pw@$      sq ~��Zݙ�q ~ q ~�9t 884t 75pw        sq ~��Zݝ�q ~ q ~�9t 884t 84pw@@�鹙�sq ~��Zݙqq ~ q ~�9t 885t 61pw        sq ~��ZݡPq ~ q ~�9t 885t 84pw@@�鹙�sq ~��Zݝ2q ~ q ~�9t 886t 61pw        sq ~��Zݥq ~ q ~�9t 886t 84pw@5oz�G�sq ~��Zݨ�q ~ q ~�9t 887t 84pw@$      sq ~��Zݬ�q ~ q ~�9t 888t 84pw@6A|CLvJsq ~��Zݬ�q ~ q ~�9t 889t 75pw        sq ~��ZݰTq ~ q ~�9t 889t 84pw@5oz�G�sq ~��W�u�q ~ q ~�9t 89t 24pw@:�+�#sq ~��W�x�q ~ q ~�9t 89t 31pw�����0Ucsq ~��WȀ�q ~ q ~�9t 89t 54pw@%��+Lsq ~��WȄ�q ~ q ~�9t 89t 67pw��ϊ��=sq ~��Wȇ�q ~ q ~�9t 89t 71pw        sq ~��Z��q ~ q ~�9t 890t 61pw        sq ~��Z��q ~ q ~�9t 890t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 891t 61pw        sq ~��Z��q ~ q ~�9t 891t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 892t 61pw        sq ~��Z�
lq ~ q ~�9t 892t 84pw@$      sq ~��Z�Nq ~ q ~�9t 893t 61pw        sq ~��Z�-q ~ q ~�9t 893t 84pw@@�鹙�sq ~��Z�
q ~ q ~�9t 894t 61pw        sq ~��Z��q ~ q ~�9t 894t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 895t 84pw@$      sq ~��Z�pq ~ q ~�9t 896t 84pw@@�鹙�sq ~��Z�Rq ~ q ~�9t 897t 61pw        sq ~��Z�1q ~ q ~�9t 897t 84pw@@�鹙�sq ~��Z�Pq ~ q ~�9t 898t 75pw        sq ~��Z� �q ~ q ~�9t 898t 84pw@5oz�G�sq ~��Z�!q ~ q ~�9t 899t 75pw        sq ~��Z�$�q ~ q ~�9t 899t 84pw@5oz�G�sq ~��W�D�q ~ q ~�9t 9t 0pw        sq ~��W�q ~ q ~�9t 9t 38pw@$      sq ~��W��q ~ q ~�9t 9t 47pw@$      sq ~��W�E;q ~ q ~�9t 9t 5pw@$      sq ~��W�ӭq ~ q ~�9t 90t 56pw@5oz�G�sq ~��W���q ~ q ~�9t 90t 74pw@5oz�G�sq ~��Z��5q ~ q ~�9t 900t 61pw        sq ~��Z�q ~ q ~�9t 900t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 901t 61pw        sq ~��Z��q ~ q ~�9t 901t 84pw@$      sq ~��Z��q ~ q ~�9t 902t 75pw        sq ~��Z�
�q ~ q ~�9t 902t 84pw@M]��%��sq ~��Z�xq ~ q ~�9t 903t 61pw        sq ~��Z�Wq ~ q ~�9t 903t 84pw@@�鹙�sq ~��Z�vq ~ q ~�9t 904t 75pw        sq ~��Z�q ~ q ~�9t 904t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 905t 61pw        sq ~��Z��q ~ q ~�9t 905t 84pw@F�U�i�sq ~��Z��q ~ q ~�9t 906t 75pw        sq ~��Z��q ~ q ~�9t 906t 84pw@F�U�i�sq ~��Z�|q ~ q ~�9t 907t 61pw        sq ~��Z�[q ~ q ~�9t 907t 84pw@@�鹙�sq ~��Z�=q ~ q ~�9t 908t 61pw        sq ~��Z�!q ~ q ~�9t 908t 84pw@@�鹙�sq ~��Z�$�q ~ q ~�9t 909t 84pw@5oz�G�sq ~��W�ڔq ~ q ~�9t 91t 61pw@$      sq ~��W���q ~ q ~�9t 91t 75pw        sq ~��W��sq ~ q ~�9t 91t 84pw@)94Go�sq ~��Z�wsq ~ q ~�9t 910t 84pw@5oz�G�sq ~��Z�sUq ~ q ~�9t 911t 61pw        sq ~��Z�{4q ~ q ~�9t 911t 84pw@@�鹙�sq ~��Z�wq ~ q ~�9t 912t 61pw        sq ~��Z�~�q ~ q ~�9t 912t 84pw@5oz�G�sq ~��Z�q ~ q ~�9t 913t 75pw        sq ~��Z肶q ~ q ~�9t 913t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 914t 75pw        sq ~��Z�wq ~ q ~�9t 914t 84pw@$      sq ~��Z�Yq ~ q ~�9t 915t 61pw        sq ~��Z�8q ~ q ~�9t 915t 84pw@5oz�G�sq ~��Z�q ~ q ~�9t 916t 61pw        sq ~��Z��q ~ q ~�9t 916t 84pw@@�鹙�sq ~��Z葺q ~ q ~�9t 917t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 918t 75pw        sq ~��Z�{q ~ q ~�9t 918t 84pw@@�鹙�sq ~��Z蕚q ~ q ~�9t 919t 75pw        sq ~��Z�<q ~ q ~�9t 919t 84pw@@�鹙�sq ~��W�Ϯq ~ q ~�9t 92t 24pw@��n@��sq ~��W��q ~ q ~�9t 92t 31pw��7��/��sq ~��W���q ~ q ~�9t 92t 53pw@$      sq ~��W���q ~ q ~�9t 92t 54pw@�^�.\sq ~��W��q ~ q ~�9t 92t 67pw���9.�Vsq ~��Z���q ~ q ~�9t 920t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 921t 75pw        sq ~��Z��q ~ q ~�9t 921t 84pw@5oz�G�sq ~��Z��Tq ~ q ~�9t 922t 84pw@5oz�G�sq ~��Z��sq ~ q ~�9t 923t 75pw        sq ~��Z��q ~ q ~�9t 923t 84pw@5oz�G�sq ~��Z��4q ~ q ~�9t 924t 75pw        sq ~��Z���q ~ q ~�9t 924t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 925t 61pw        sq ~��Z���q ~ q ~�9t 925t 84pw@5oz�G�sq ~��Z��yq ~ q ~�9t 926t 61pw        sq ~��Z�Xq ~ q ~�9t 926t 84pw@5oz�G�sq ~��Z�q ~ q ~�9t 927t 84pw@@�鹙�sq ~��Z�8q ~ q ~�9t 928t 75pw        sq ~��Z�	�q ~ q ~�9t 928t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 929t 61pw        sq ~��Z��q ~ q ~�9t 929t 84pw@@�鹙�sq ~��W�`q ~ q ~�9t 93t 1pw@&n��:ssq ~��W��5q ~ q ~�9t 93t 62pw        sq ~��Z�\�q ~ q ~�9t 930t 75pw        sq ~��Z�`1q ~ q ~�9t 930t 84pw@$      sq ~��Z�\q ~ q ~�9t 931t 61pw        sq ~��Z�c�q ~ q ~�9t 931t 84pw@$      sq ~��Z�_�q ~ q ~�9t 932t 61pw        sq ~��Z�g�q ~ q ~�9t 932t 84pw@5oz�G�sq ~��Z�c�q ~ q ~�9t 933t 61pw        sq ~��Z�ktq ~ q ~�9t 933t 84pw@@�鹙�sq ~��Z�k�q ~ q ~�9t 934t 75pw        sq ~��Z�o5q ~ q ~�9t 934t 84pw@5oz�G�sq ~��Z�kq ~ q ~�9t 935t 61pw        sq ~��Z�r�q ~ q ~�9t 935t 84pw@5oz�G�sq ~��Z�n�q ~ q ~�9t 936t 61pw        sq ~��Z�v�q ~ q ~�9t 936t 84pw@5oz�G�sq ~��Z�r�q ~ q ~�9t 937t 61pw        sq ~��Z�zxq ~ q ~�9t 937t 84pw@$      sq ~��Z�~9q ~ q ~�9t 938t 84pw@@�鹙�sq ~��Z�~Xq ~ q ~�9t 939t 75pw        sq ~��Z��q ~ q ~�9t 939t 84pw@@�鹙�sq ~��W�׍q ~ q ~�9t 94t 27pw@!^ƪT��sq ~��Z�̱q ~ q ~�9t 940t 61pw        sq ~��Z�Ԑq ~ q ~�9t 940t 84pw@$      sq ~��Z��Qq ~ q ~�9t 941t 84pw@$#�a�
sq ~��Z��3q ~ q ~�9t 942t 61pw        sq ~��Z��q ~ q ~�9t 942t 84pw@F�U�i�sq ~��Z��1q ~ q ~�9t 943t 75pw        sq ~��Z���q ~ q ~�9t 943t 84pw@@�鹙�sq ~��Z�۵q ~ q ~�9t 944t 61pw        sq ~��Z��q ~ q ~�9t 944t 84pw@@�鹙�sq ~��Z��Uq ~ q ~�9t 945t 84pw@@�鹙�sq ~��Z��7q ~ q ~�9t 946t 61pw        sq ~��Z��q ~ q ~�9t 946t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 947t 61pw        sq ~��Z���q ~ q ~�9t 947t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 948t 75pw        sq ~��Z��q ~ q ~�9t 948t 84pw@$      sq ~��Z��Yq ~ q ~�9t 949t 84pw@$      sq ~��W��Nq ~ q ~�9t 95t 27pw?�3�_�sq ~��Z�H�q ~ q ~�9t 950t 84pw@5oz�G�sq ~��Z�Iq ~ q ~�9t 951t 75pw        sq ~��Z�L�q ~ q ~�9t 951t 84pw@$      sq ~��Z�H�q ~ q ~�9t 952t 61pw        sq ~��Z�Pqq ~ q ~�9t 952t 84pw@$      sq ~��Z�P�q ~ q ~�9t 953t 75pw        sq ~��Z�T2q ~ q ~�9t 953t 84pw@@�鹙�sq ~��Z�TQq ~ q ~�9t 954t 75pw        sq ~��Z�W�q ~ q ~�9t 954t 84pw@5oz�G�sq ~��Z�Xq ~ q ~�9t 955t 75pw        sq ~��Z�[�q ~ q ~�9t 955t 84pw@@�鹙�sq ~��Z�W�q ~ q ~�9t 956t 61pw        sq ~��Z�_uq ~ q ~�9t 956t 84pw@@�鹙�sq ~��Z�_�q ~ q ~�9t 957t 75pw        sq ~��Z�c6q ~ q ~�9t 957t 84pw@@�鹙�sq ~��Z�_q ~ q ~�9t 958t 61pw        sq ~��Z�f�q ~ q ~�9t 958t 84pw@5oz�G�sq ~��Z�b�q ~ q ~�9t 959t 61pw        sq ~��Z�j�q ~ q ~�9t 959t 84pw@@�鹙�sq ~��W��q ~ q ~�9t 96t 27pw@%��*��sq ~��W��:q ~ q ~�9t 96t 60pw        sq ~��W��2q ~ q ~�9t 96t 68pw��T~ȯ%sq ~��Z�oq ~ q ~�9t 960t 61pw        sq ~��Z�Nq ~ q ~�9t 960t 84pw@F�U�i�sq ~��Z�0q ~ q ~�9t 961t 61pw        sq ~��Z��q ~ q ~�9t 961t 84pw@$      sq ~��Z��q ~ q ~�9t 962t 61pw        sq ~��Z���q ~ q ~�9t 962t 84pw@5oz�G�sq ~��Z���q ~ q ~�9t 963t 61pw        sq ~��Z�ȑq ~ q ~�9t 963t 84pw@F�U�i�sq ~��Z��sq ~ q ~�9t 964t 61pw        sq ~��Z��Rq ~ q ~�9t 964t 84pw@@�鹙�sq ~��Z��4q ~ q ~�9t 965t 61pw        sq ~��Z��q ~ q ~�9t 965t 84pw@@�鹙�sq ~��Z���q ~ q ~�9t 966t 84pw@@�鹙�sq ~��Z�϶q ~ q ~�9t 967t 61pw        sq ~��Z�וq ~ q ~�9t 967t 84pw@5oz�G�sq ~��Z�״q ~ q ~�9t 968t 75pw        sq ~��Z��Vq ~ q ~�9t 968t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 969t 84pw@$      sq ~��W���q ~ q ~�9t 97t 77pw@@�鹙�sq ~��Z�.q ~ q ~�9t 970t 75pw        sq ~��Z�1�q ~ q ~�9t 970t 84pw@$      sq ~��Z�1�q ~ q ~�9t 971t 75pw        sq ~��Z�5nq ~ q ~�9t 971t 84pw@5oz�G�sq ~��Z�5�q ~ q ~�9t 972t 75pw        sq ~��Z�9/q ~ q ~�9t 972t 84pw@$      sq ~��Z�9Nq ~ q ~�9t 973t 75pw        sq ~��Z�<�q ~ q ~�9t 973t 84pw@5oz�G�sq ~��Z�=q ~ q ~�9t 974t 75pw        sq ~��Z�@�q ~ q ~�9t 974t 84pw@5oz�G�sq ~��Z�@�q ~ q ~�9t 975t 75pw        sq ~��Z�Drq ~ q ~�9t 975t 84pw@5oz�G�sq ~��Z�D�q ~ q ~�9t 976t 75pw        sq ~��Z�H3q ~ q ~�9t 976t 84pw@$      sq ~��Z�HRq ~ q ~�9t 977t 75pw        sq ~��Z�K�q ~ q ~�9t 977t 84pw@5oz�G�sq ~��Z�Lq ~ q ~�9t 978t 75pw        sq ~��Z�O�q ~ q ~�9t 978t 84pw@@�鹙�sq ~��Z�Svq ~ q ~�9t 979t 84pw@5oz�G�sq ~��W��uq ~ q ~�9t 98t 78pw@:����sq ~��Z�-q ~ q ~�9t 980t 61pw        sq ~��Z�q ~ q ~�9t 980t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 981t 84pw@5oz�G�sq ~��Z��q ~ q ~�9t 982t 75pw        sq ~��Z뭎q ~ q ~�9t 982t 84pw@$      sq ~��Z뭭q ~ q ~�9t 983t 75pw        sq ~��Z�Oq ~ q ~�9t 983t 84pw@$      sq ~��Z�nq ~ q ~�9t 984t 75pw        sq ~��Z�q ~ q ~�9t 984t 84pw@$      sq ~��Z�/q ~ q ~�9t 985t 75pw        sq ~��Z��q ~ q ~�9t 985t 84pw@5oz�G�sq ~��Z봳q ~ q ~�9t 986t 61pw        sq ~��Z뼒q ~ q ~�9t 986t 84pw@$      sq ~��Z��Sq ~ q ~�9t 987t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 988t 84pw@$      sq ~��Z��q ~ q ~�9t 989t 61pw        sq ~��Z���q ~ q ~�9t 989t 84pw@5oz�G�sq ~��W��vq ~ q ~�9t 99t 56pw@/^�K,��sq ~��W���q ~ q ~�9t 99t 74pw@$�
υ�bsq ~��Z�kq ~ q ~�9t 990t 84pw@@�鹙�sq ~��Z�,q ~ q ~�9t 991t 84pw@5oz�G�sq ~��Z�!�q ~ q ~�9t 992t 84pw@@�鹙�sq ~��Z��q ~ q ~�9t 993t 61pw        sq ~��Z�%�q ~ q ~�9t 993t 84pw@5oz�G�sq ~��Z�!�q ~ q ~�9t 994t 61pw        sq ~��Z�)oq ~ q ~�9t 994t 84pw@@�鹙�sq ~��Z�-0q ~ q ~�9t 995t 84pw@@�鹙�sq ~��Z�0�q ~ q ~�9t 996t 84pw@@�鹙�sq ~��Z�4�q ~ q ~�9t 997t 84pw@5oz�G�sq ~��Z�0�q ~ q ~�9t 998t 61pw        sq ~��Z�8sq ~ q ~�9t 998t 84pw@$      sq ~��Z�4Uq ~ q ~�9t 999t 61pw        sq ~��Z�<4q ~ q ~�9t 999t 84pw@@�鹙�q ~��w?�      sq ~��e��q ~ t TMPt 0ppw��g4���sq ~��e���q ~ q ~�mt 1ppw?��a!!�sq ~��e�A>q ~ q ~�mt 10ppw��u����sq ~��e�D�q ~ q ~�mt 11ppw        sq ~��e�H�q ~ q ~�mt 12ppw@ %b���?sq ~��e�L�q ~ q ~�mt 13ppw?��FY�,sq ~��e�PBq ~ q ~�mt 14ppw@

|sq ~��e�Tq ~ q ~�mt 15ppw��-��)u�sq ~��e�W�q ~ q ~�mt 16ppw?�;�;Аsq ~��e�[�q ~ q ~�mt 17ppw?�3�,�U�sq ~��e�_Fq ~ q ~�mt 18ppw?��#���sq ~��e�cq ~ q ~�mt 19ppw?�M?�sq ~��e��q ~ q ~�mt 2ppw?���[gVsq ~��eص�q ~ q ~�mt 20ppw        sq ~��eع^q ~ q ~�mt 21ppw?�
�7��&sq ~��eؽq ~ q ~�mt 22ppw@��_8P�sq ~��e���q ~ q ~�mt 23ppw?�JЏ�sq ~��e�ġq ~ q ~�mt 24ppw?��4&���sq ~��e��bq ~ q ~�mt 25ppw?�2�.{��sq ~��e��#q ~ q ~�mt 26ppw?ޑ�����sq ~��e���q ~ q ~�mt 27ppw@��5?�sq ~��e�ӥq ~ q ~�mt 28ppw?��1��Wsq ~��e��fq ~ q ~�mt 29ppw��m�"��sq ~��e�Rq ~ q ~�mt 3ppw���}߉�sq ~��e�)�q ~ q ~�mt 30ppw?�JĽa�sq ~��e�-�q ~ q ~�mt 31ppw��._�@�sq ~��e�1~q ~ q ~�mt 32ppw?u��9ȁsq ~��e�5?q ~ q ~�mt 33ppw��Ht�k�sq ~��e�9 q ~ q ~�mt 34ppw        sq ~��e�<�q ~ q ~�mt 35ppw��;����sq ~��e�@�q ~ q ~�mt 36ppw��4�~ûsq ~��e�DCq ~ q ~�mt 37ppw����@��sq ~��e�Hq ~ q ~�mt 38ppw@�%�8sq ~��e�K�q ~ q ~�mt 39ppw?�!��I�Dsq ~��e�
q ~ q ~�mt 4ppw���ˋY��sq ~��eٞ[q ~ q ~�mt 40ppw?�G�^��lsq ~��e٢q ~ q ~�mt 41ppw?�7|�g�sq ~��e٥�q ~ q ~�mt 42ppw        sq ~��e٩�q ~ q ~�mt 43ppw��+,3�vsq ~��e٭_q ~ q ~�mt 44ppw?�_'��4�sq ~��eٱ q ~ q ~�mt 45ppw?���6sq ~��eٴ�q ~ q ~�mt 46ppw?��2��sq ~��eٸ�q ~ q ~�mt 47ppw?�D���<sq ~��eټcq ~ q ~�mt 48ppw?��d�$Jsq ~��e��$q ~ q ~�mt 49ppw?�4_ ��Gsq ~��e��q ~ q ~�mt 5ppw���J�cP�sq ~��e��q ~ q ~�mt 50ppw?���&�sq ~��e�{q ~ q ~�mt 51ppw?�H-d�>sq ~��e�<q ~ q ~�mt 52ppw��;����sq ~��e��q ~ q ~�mt 53ppw?�T�ErYsq ~��e�!�q ~ q ~�mt 54ppw?�
�2�h�sq ~��e�%q ~ q ~�mt 55ppw        sq ~��e�)@q ~ q ~�mt 56ppw?��2l��sq ~��e�-q ~ q ~�mt 57ppw?�P%=�sq ~��e�0�q ~ q ~�mt 58ppw        sq ~��e�4�q ~ q ~�mt 59ppw��ͤ[.esq ~��e��q ~ q ~�mt 6ppw@Q
��sq ~��eڇq ~ q ~�mt 60ppw?�g
��?sq ~��eڊ�q ~ q ~�mt 61ppw����a7 }sq ~��eڎ�q ~ q ~�mt 62ppw        sq ~��eڒ\q ~ q ~�mt 63ppw��J�
s��sq ~��eږq ~ q ~�mt 64ppw?��d�$Jsq ~��eڙ�q ~ q ~�mt 65ppw?������&sq ~��eڝ�q ~ q ~�mt 66ppw        sq ~��eڡ`q ~ q ~�mt 67ppw��z7H�sq ~��eڥ!q ~ q ~�mt 68ppw?�ݽ�~�@sq ~��eڨ�q ~ q ~�mt 69ppw        sq ~��e�Vq ~ q ~�mt 7ppw����!��sq ~��e��xq ~ q ~�mt 70ppw        sq ~��e��9q ~ q ~�mt 71ppw        sq ~��e��q ~ q ~�mt 72ppw��#�,��Jsq ~��e��q ~ q ~�mt 73ppw?�v���.sq ~��e�
|q ~ q ~�mt 74ppw?���m�2�sq ~��e�=q ~ q ~�mt 75ppw        sq ~��e��q ~ q ~�mt 76ppw        sq ~��e��q ~ q ~�mt 77ppw        sq ~��e��q ~ q ~�mt 78ppw?�4|^_I=sq ~��e�Aq ~ q ~�mt 79ppw        sq ~��e�q ~ q ~�mt 8ppw?����H�fsq ~��e�o�q ~ q ~�mt 80ppw?�4_ ��Gsq ~��e�s�q ~ q ~�mt 81ppw        sq ~��e�wYq ~ q ~�mt 82ppw?����sq ~��e�{q ~ q ~�mt 83ppw?�4_ ��Gsq ~��e�~�q ~ q ~�mt 84ppw@��2�Zsq ~��e��q ~ q ~�mt 9ppw?ᣊ/uq ~��w?�      sq ~��{H�q ~ t XEMEt 0ppw@$      sq ~��{H��q ~ q ~�t 1ppw@$      sq ~��{^�0q ~ q ~�t 10ppw@%���}B�sq ~��~��q ~ q ~�t 100ppw@.�B���)sq ~��ѠXpq ~ q ~�t 1000ppw@$      sq ~��Ѡ\1q ~ q ~�t 1001ppw@$      sq ~��Ѡ_�q ~ q ~�t 1002ppw@$      sq ~��Ѡc�q ~ q ~�t 1003ppw@$      sq ~��Ѡgtq ~ q ~�t 1004ppw@$      sq ~��Ѡk5q ~ q ~�t 1005ppw@$      sq ~��Ѡn�q ~ q ~�t 1006ppw@$      sq ~��Ѡr�q ~ q ~�t 1007ppw@$      sq ~��Ѡvxq ~ q ~�t 1008ppw@$      sq ~��Ѡz9q ~ q ~�t 1009ppw@$      sq ~��~�Cq ~ q ~�t 101ppw@$      sq ~��Ѡ��q ~ q ~�t 1010ppw@$      sq ~��ѠАq ~ q ~�t 1011ppw@$      sq ~��Ѡ�Qq ~ q ~�t 1012ppw@$      sq ~��Ѡ�q ~ q ~�t 1013ppw@$      sq ~��Ѡ��q ~ q ~�t 1014ppw@$      sq ~��Ѡߔq ~ q ~�t 1015ppw@$      sq ~��Ѡ�Uq ~ q ~�t 1016ppw@$      sq ~��Ѡ�q ~ q ~�t 1017ppw@$      sq ~��Ѡ��q ~ q ~�t 1018ppw@$      sq ~��Ѡ�q ~ q ~�t 1019ppw@$      sq ~��~q ~ q ~�t 102ppw@$      sq ~��ѡA.q ~ q ~�t 1020ppw@$      sq ~��ѡD�q ~ q ~�t 1021ppw@$      sq ~��ѡH�q ~ q ~�t 1022ppw@$      sq ~��ѡLqq ~ q ~�t 1023ppw@$      sq ~��ѡP2q ~ q ~�t 1024ppw@$      sq ~��ѡS�q ~ q ~�t 1025ppw@$      sq ~��ѡW�q ~ q ~�t 1026ppw@$      sq ~��ѡ[uq ~ q ~�t 1027ppw@$      sq ~��ѡ_6q ~ q ~�t 1028ppw@$      sq ~��ѡb�q ~ q ~�t 1029ppw@$      sq ~��~�q ~ q ~�t 103ppw@$      sq ~��ѡ��q ~ q ~�t 1030ppw@$      sq ~��ѡ�Nq ~ q ~�t 1031ppw@$      sq ~��ѡ�q ~ q ~�t 1032ppw@$      sq ~��ѡ��q ~ q ~�t 1033ppw@$      sq ~��ѡđq ~ q ~�t 1034ppw@$      sq ~��ѡ�Rq ~ q ~�t 1035ppw@$      sq ~��ѡ�q ~ q ~�t 1036ppw@$      sq ~��ѡ��q ~ q ~�t 1037ppw@$      sq ~��ѡӕq ~ q ~�t 1038ppw@$      sq ~��ѡ�Vq ~ q ~�t 1039ppw@$      sq ~��~�q ~ q ~�t 104ppw@$      sq ~��Ѣ)�q ~ q ~�t 1040ppw@$      sq ~��Ѣ-�q ~ q ~�t 1041ppw@$      sq ~��Ѣ1nq ~ q ~�t 1042ppw@$      sq ~��Ѣ5/q ~ q ~�t 1043ppw@$      sq ~��Ѣ8�q ~ q ~�t 1044ppw@$      sq ~��Ѣ<�q ~ q ~�t 1045ppw@$      sq ~��Ѣ@rq ~ q ~�t 1046ppw@$      sq ~��ѢD3q ~ q ~�t 1047ppw@$      sq ~��ѢG�q ~ q ~�t 1048ppw@$      sq ~��ѢK�q ~ q ~�t 1049ppw@$      sq ~��~Gq ~ q ~�t 105ppw@$      sq ~��Ѣ�Kq ~ q ~�t 1050ppw@$      sq ~��Ѣ�q ~ q ~�t 1051ppw@$      sq ~��Ѣ��q ~ q ~�t 1052ppw@$      sq ~��Ѣ��q ~ q ~�t 1053ppw@$      sq ~��Ѣ�Oq ~ q ~�t 1054ppw@$      sq ~��Ѣ�q ~ q ~�t 1055ppw@$      sq ~��Ѣ��q ~ q ~�t 1056ppw@$      sq ~��Ѣ��q ~ q ~�t 1057ppw@$      sq ~��Ѣ�Sq ~ q ~�t 1058ppw@$      sq ~��Ѣ�q ~ q ~�t 1059ppw@$      sq ~��~q ~ q ~�t 106ppw@$      sq ~��ѣ�q ~ q ~�t 1060ppw@$      sq ~��ѣkq ~ q ~�t 1061ppw@$      sq ~��ѣ,q ~ q ~�t 1062ppw@$      sq ~��ѣ�q ~ q ~�t 1063ppw@$      sq ~��ѣ!�q ~ q ~�t 1064ppw@$      sq ~��ѣ%oq ~ q ~�t 1065ppw@$      sq ~��ѣ)0q ~ q ~�t 1066ppw@$      sq ~��ѣ,�q ~ q ~�t 1067ppw@#�K`�Esq ~��ѣ0�q ~ q ~�t 1068ppw@$      sq ~��ѣ4sq ~ q ~�t 1069ppw@$      sq ~��~�q ~ q ~�t 107ppw@$      sq ~��ѣ�	q ~ q ~�t 1070ppw@$      sq ~��ѣ��q ~ q ~�t 1071ppw@$      sq ~��ѣ��q ~ q ~�t 1072ppw@$      sq ~��ѣ�Lq ~ q ~�t 1073ppw@$      sq ~��ѣ�q ~ q ~�t 1074ppw@$      sq ~��ѣ��q ~ q ~�t 1075ppw@$      sq ~��ѣ��q ~ q ~�t 1076ppw@$      sq ~��ѣ�Pq ~ q ~�t 1077ppw@$      sq ~��ѣ�q ~ q ~�t 1078ppw@$      sq ~��ѣ��q ~ q ~�t 1079ppw@$      sq ~��~�q ~ q ~�t 108ppw@$      sq ~��ѣ�hq ~ q ~�t 1080ppw@$      sq ~��ѣ�)q ~ q ~�t 1081ppw@$      sq ~��Ѥ�q ~ q ~�t 1082ppw@$      sq ~��Ѥ�q ~ q ~�t 1083ppw@$      sq ~��Ѥ
lq ~ q ~�t 1084ppw@$      sq ~��Ѥ-q ~ q ~�t 1085ppw@$      sq ~��Ѥ�q ~ q ~�t 1086ppw@$      sq ~��Ѥ�q ~ q ~�t 1087ppw@$      sq ~��Ѥpq ~ q ~�t 1088ppw@$      sq ~��Ѥ1q ~ q ~�t 1089ppw@$      sq ~��~Kq ~ q ~�t 109ppw@$      sq ~��Ѥo�q ~ q ~�t 1090ppw@$      sq ~��Ѥs�q ~ q ~�t 1091ppw@$      sq ~��ѤwIq ~ q ~�t 1092ppw@$      sq ~��Ѥ{
q ~ q ~�t 1093ppw@$      sq ~��Ѥ~�q ~ q ~�t 1094ppw@$      sq ~��Ѥ��q ~ q ~�t 1095ppw@$      sq ~��Ѥ�Mq ~ q ~�t 1096ppw@$      sq ~��Ѥ�q ~ q ~�t 1097ppw@$      sq ~��Ѥ��q ~ q ~�t 1098ppw@$      sq ~��Ѥ��q ~ q ~�t 1099ppw@$      sq ~��{^��q ~ q ~�t 11ppw@/��ܷsq ~��~m�q ~ q ~�t 110ppw@$      sq ~��Ѯo�q ~ q ~�t 1100ppw@$      sq ~��Ѯs�q ~ q ~�t 1101ppw@$      sq ~��Ѯwsq ~ q ~�t 1102ppw@$      sq ~��Ѯ{4q ~ q ~�t 1103ppw@$      sq ~��Ѯ~�q ~ q ~�t 1104ppw@$      sq ~��Ѯ��q ~ q ~�t 1105ppw@#�ϗ�X�sq ~��Ѯ�wq ~ q ~�t 1106ppw@$      sq ~��Ѯ�8q ~ q ~�t 1107ppw@$      sq ~��Ѯ��q ~ q ~�t 1108ppw@$      sq ~��Ѯ��q ~ q ~�t 1109ppw@$      sq ~��~q�q ~ q ~�t 111ppw@$      sq ~��Ѯ�Pq ~ q ~�t 1110ppw@$      sq ~��Ѯ�q ~ q ~�t 1111ppw@$      sq ~��Ѯ��q ~ q ~�t 1112ppw@$      sq ~��Ѯ�q ~ q ~�t 1113ppw@$      sq ~��Ѯ�Tq ~ q ~�t 1114ppw@$      sq ~��Ѯ�q ~ q ~�t 1115ppw@$      sq ~��Ѯ��q ~ q ~�t 1116ppw@#��W�6sq ~��Ѯ��q ~ q ~�t 1117ppw@$      sq ~��ѯXq ~ q ~�t 1118ppw@$      sq ~��ѯq ~ q ~�t 1119ppw@$      sq ~��~ucq ~ q ~�t 112ppw@$      sq ~��ѯX�q ~ q ~�t 1120ppw@$      sq ~��ѯ\pq ~ q ~�t 1121ppw@$      sq ~��ѯ`1q ~ q ~�t 1122ppw@$      sq ~��ѯc�q ~ q ~�t 1123ppw@'���jsq ~��ѯg�q ~ q ~�t 1124ppw@$      sq ~��ѯktq ~ q ~�t 1125ppw@$      sq ~��ѯo5q ~ q ~�t 1126ppw@$      sq ~��ѯr�q ~ q ~�t 1127ppw@$      sq ~��ѯv�q ~ q ~�t 1128ppw@$      sq ~��ѯzxq ~ q ~�t 1129ppw@$      sq ~��~y$q ~ q ~�t 113ppw@$      sq ~��ѯ�q ~ q ~�t 1130ppw@$��G74sq ~��ѯ��q ~ q ~�t 1131ppw@%�����ksq ~��ѯԐq ~ q ~�t 1132ppw@$      sq ~��ѯ�Qq ~ q ~�t 1133ppw@$      sq ~��ѯ�q ~ q ~�t 1134ppw@$      sq ~��ѯ��q ~ q ~�t 1135ppw@$      sq ~��ѯ�q ~ q ~�t 1136ppw@$      sq ~��ѯ�Uq ~ q ~�t 1137ppw@$      sq ~��ѯ�q ~ q ~�t 1138ppw@$      sq ~��ѯ��q ~ q ~�t 1139ppw@$      sq ~��~|�q ~ q ~�t 114ppw@%�1T�a[sq ~��ѰAmq ~ q ~�t 1140ppw@$      sq ~��ѰE.q ~ q ~�t 1141ppw@$      sq ~��ѰH�q ~ q ~�t 1142ppw@$      sq ~��ѰL�q ~ q ~�t 1143ppw@$      sq ~��ѰPqq ~ q ~�t 1144ppw@$      sq ~��ѰT2q ~ q ~�t 1145ppw@$      sq ~��ѰW�q ~ q ~�t 1146ppw@$      sq ~��Ѱ[�q ~ q ~�t 1147ppw@$      sq ~��Ѱ_uq ~ q ~�t 1148ppw@$      sq ~��Ѱc6q ~ q ~�t 1149ppw@$      sq ~��~��q ~ q ~�t 115ppw@$      sq ~��Ѱ��q ~ q ~�t 1150ppw@$      sq ~��Ѱ��q ~ q ~�t 1151ppw@$      sq ~��Ѱ�Nq ~ q ~�t 1152ppw@$      sq ~��Ѱ�q ~ q ~�t 1153ppw@$      sq ~��Ѱ��q ~ q ~�t 1154ppw@$      sq ~��Ѱȑq ~ q ~�t 1155ppw@$      sq ~��Ѱ�Rq ~ q ~�t 1156ppw@$      sq ~��Ѱ�q ~ q ~�t 1157ppw@$      sq ~��Ѱ��q ~ q ~�t 1158ppw@$      sq ~��Ѱוq ~ q ~�t 1159ppw@$      sq ~��~�gq ~ q ~�t 116ppw@$      sq ~��ѱ*+q ~ q ~�t 1160ppw@"D�^���sq ~��ѱ-�q ~ q ~�t 1161ppw@$      sq ~��ѱ1�q ~ q ~�t 1162ppw@$      sq ~��ѱ5nq ~ q ~�t 1163ppw@$      sq ~��ѱ9/q ~ q ~�t 1164ppw@$      sq ~��ѱ<�q ~ q ~�t 1165ppw@$      sq ~��ѱ@�q ~ q ~�t 1166ppw@$      sq ~��ѱDrq ~ q ~�t 1167ppw@$      sq ~��ѱH3q ~ q ~�t 1168ppw@$      sq ~��ѱK�q ~ q ~�t 1169ppw@$      sq ~��~�(q ~ q ~�t 117ppw@$      sq ~��ѱ��q ~ q ~�t 1170ppw@$      sq ~��ѱ�Kq ~ q ~�t 1171ppw@$      sq ~��ѱ�q ~ q ~�t 1172ppw@$      sq ~��ѱ��q ~ q ~�t 1173ppw@$      sq ~��ѱ��q ~ q ~�t 1174ppw@$      sq ~��ѱ�Oq ~ q ~�t 1175ppw@$      sq ~��ѱ�q ~ q ~�t 1176ppw@$      sq ~��ѱ��q ~ q ~�t 1177ppw@$      sq ~��ѱ��q ~ q ~�t 1178ppw@$      sq ~��ѱ�Sq ~ q ~�t 1179ppw@$      sq ~��~��q ~ q ~�t 118ppw@$      sq ~��Ѳ�q ~ q ~�t 1180ppw@$      sq ~��Ѳ�q ~ q ~�t 1181ppw@$      sq ~��Ѳkq ~ q ~�t 1182ppw@$      sq ~��Ѳ,q ~ q ~�t 1183ppw@$      sq ~��Ѳ!�q ~ q ~�t 1184ppw@$      sq ~��Ѳ%�q ~ q ~�t 1185ppw@$      sq ~��Ѳ)oq ~ q ~�t 1186ppw@$      sq ~��Ѳ-0q ~ q ~�t 1187ppw@$      sq ~��Ѳ0�q ~ q ~�t 1188ppw@$      sq ~��Ѳ4�q ~ q ~�t 1189ppw@$      sq ~��~��q ~ q ~�t 119ppw@$      sq ~��Ѳ�Hq ~ q ~�t 1190ppw@$      sq ~��Ѳ�	q ~ q ~�t 1191ppw@$      sq ~��Ѳ��q ~ q ~�t 1192ppw@$      sq ~��Ѳ��q ~ q ~�t 1193ppw@$      sq ~��Ѳ�Lq ~ q ~�t 1194ppw@$      sq ~��Ѳ�q ~ q ~�t 1195ppw@$      sq ~��Ѳ��q ~ q ~�t 1196ppw@'�p��j�sq ~��Ѳ��q ~ q ~�t 1197ppw@$      sq ~��Ѳ�Pq ~ q ~�t 1198ppw@$      sq ~��Ѳ�q ~ q ~�t 1199ppw@$      sq ~��{^��q ~ q ~�t 12ppw@$      sq ~��~�@q ~ q ~�t 120ppw@$      sq ~��Ѽ�rq ~ q ~�t 1200ppw@$      sq ~��Ѽ�3q ~ q ~�t 1201ppw@$      sq ~��Ѽ��q ~ q ~�t 1202ppw@$      sq ~��Ѽ��q ~ q ~�t 1203ppw@$      sq ~��Ѽ�vq ~ q ~�t 1204ppw@$      sq ~��Ѽ�7q ~ q ~�t 1205ppw@$      sq ~��Ѽ��q ~ q ~�t 1206ppw@$      sq ~��Ѽ��q ~ q ~�t 1207ppw@$      sq ~��Ѽ�zq ~ q ~�t 1208ppw@$      sq ~��Ѽ�;q ~ q ~�t 1209ppw@$      sq ~��~�q ~ q ~�t 121ppw@$      sq ~��Ѽ��q ~ q ~�t 1210ppw@$      sq ~��Ѽ��q ~ q ~�t 1211ppw@$      sq ~��ѽSq ~ q ~�t 1212ppw@$      sq ~��ѽq ~ q ~�t 1213ppw@$      sq ~��ѽ
�q ~ q ~�t 1214ppw@$      sq ~��ѽ�q ~ q ~�t 1215ppw@$      sq ~��ѽWq ~ q ~�t 1216ppw@$      sq ~��ѽq ~ q ~�t 1217ppw@$      sq ~��ѽ�q ~ q ~�t 1218ppw@$      sq ~��ѽ�q ~ q ~�t 1219ppw@$      sq ~��~��q ~ q ~�t 122ppw@$      sq ~��ѽp0q ~ q ~�t 1220ppw@$      sq ~��ѽs�q ~ q ~�t 1221ppw@$      sq ~��ѽw�q ~ q ~�t 1222ppw@$      sq ~��ѽ{sq ~ q ~�t 1223ppw@$      sq ~��ѽ4q ~ q ~�t 1224ppw@$      sq ~��ѽ��q ~ q ~�t 1225ppw@$      sq ~��ѽ��q ~ q ~�t 1226ppw@$      sq ~��ѽ�wq ~ q ~�t 1227ppw@$      sq ~��ѽ�8q ~ q ~�t 1228ppw@$      sq ~��ѽ��q ~ q ~�t 1229ppw@$      sq ~��~�q ~ q ~�t 123ppw@$      sq ~��ѽ�q ~ q ~�t 1230ppw@$      sq ~��ѽ�Pq ~ q ~�t 1231ppw@$      sq ~��ѽ�q ~ q ~�t 1232ppw@$      sq ~��ѽ��q ~ q ~�t 1233ppw@$      sq ~��ѽ�q ~ q ~�t 1234ppw@$      sq ~��ѽ�Tq ~ q ~�t 1235ppw@$      sq ~��ѽ�q ~ q ~�t 1236ppw@$      sq ~��ѽ��q ~ q ~�t 1237ppw@$      sq ~��Ѿ�q ~ q ~�t 1238ppw@$      sq ~��ѾXq ~ q ~�t 1239ppw@$      sq ~��~�Dq ~ q ~�t 124ppw@$      sq ~��ѾX�q ~ q ~�t 1240ppw@$      sq ~��Ѿ\�q ~ q ~�t 1241ppw@#�׭�Bsq ~��Ѿ`pq ~ q ~�t 1242ppw@$      sq ~��Ѿd1q ~ q ~�t 1243ppw@$      sq ~��Ѿg�q ~ q ~�t 1244ppw@$      sq ~��Ѿk�q ~ q ~�t 1245ppw@$      sq ~��Ѿotq ~ q ~�t 1246ppw@$      sq ~��Ѿs5q ~ q ~�t 1247ppw@$      sq ~��Ѿv�q ~ q ~�t 1248ppw@$      sq ~��Ѿz�q ~ q ~�t 1249ppw@$      sq ~��~�q ~ q ~�t 125ppw@$      sq ~��Ѿ�Mq ~ q ~�t 1250ppw@$      sq ~��Ѿ�q ~ q ~�t 1251ppw@$      sq ~��Ѿ��q ~ q ~�t 1252ppw@$      sq ~��Ѿؐq ~ q ~�t 1253ppw@$      sq ~��Ѿ�Qq ~ q ~�t 1254ppw@$      sq ~��Ѿ�q ~ q ~�t 1255ppw@$      sq ~��Ѿ��q ~ q ~�t 1256ppw@$      sq ~��Ѿ�q ~ q ~�t 1257ppw@#3���sq ~��Ѿ�Uq ~ q ~�t 1258ppw@#�����Jsq ~��Ѿ�q ~ q ~�t 1259ppw@$      sq ~��~��q ~ q ~�t 126ppw@$      sq ~��ѿA�q ~ q ~�t 1260ppw@$      sq ~��ѿEmq ~ q ~�t 1261ppw@$      sq ~��ѿI.q ~ q ~�t 1262ppw@$      sq ~��ѿL�q ~ q ~�t 1263ppw@$      sq ~��ѿP�q ~ q ~�t 1264ppw@$      sq ~��ѿTqq ~ q ~�t 1265ppw@$      sq ~��ѿX2q ~ q ~�t 1266ppw@$      sq ~��ѿ[�q ~ q ~�t 1267ppw@$      sq ~��ѿ_�q ~ q ~�t 1268ppw@$      sq ~��ѿcuq ~ q ~�t 1269ppw@$      sq ~��~��q ~ q ~�t 127ppw@$      sq ~��ѿ�q ~ q ~�t 1270ppw@$      sq ~��ѿ��q ~ q ~�t 1271ppw@$      sq ~��ѿ��q ~ q ~�t 1272ppw@$      sq ~��ѿ�Nq ~ q ~�t 1273ppw@$      sq ~��ѿ�q ~ q ~�t 1274ppw@$      sq ~��ѿ��q ~ q ~�t 1275ppw@$      sq ~��ѿ̑q ~ q ~�t 1276ppw@$      sq ~��ѿ�Rq ~ q ~�t 1277ppw@$      sq ~��ѿ�q ~ q ~�t 1278ppw@+�,W8�*sq ~��ѿ��q ~ q ~�t 1279ppw@$      sq ~��~ Hq ~ q ~�t 128ppw@$      sq ~����*jq ~ q ~�t 1280ppw@$      sq ~����.+q ~ q ~�t 1281ppw@$      sq ~����1�q ~ q ~�t 1282ppw@$      sq ~����5�q ~ q ~�t 1283ppw@$      sq ~����9nq ~ q ~�t 1284ppw@$      sq ~����=/q ~ q ~�t 1285ppw@$      sq ~����@�q ~ q ~�t 1286ppw@$      sq ~����D�q ~ q ~�t 1287ppw@$      sq ~����Hrq ~ q ~�t 1288ppw@$      sq ~����L3q ~ q ~�t 1289ppw@$      sq ~��~	q ~ q ~�t 129ppw@$      sq ~������q ~ q ~�t 1290ppw@$      sq ~������q ~ q ~�t 1291ppw@$      sq ~�����Kq ~ q ~�t 1292ppw@$      sq ~�����q ~ q ~�t 1293ppw@$      sq ~������q ~ q ~�t 1294ppw@$      sq ~������q ~ q ~�t 1295ppw@$      sq ~�����Oq ~ q ~�t 1296ppw@$      sq ~�����q ~ q ~�t 1297ppw@$      sq ~������q ~ q ~�t 1298ppw@$      sq ~������q ~ q ~�t 1299ppw@$      sq ~��{^�sq ~ q ~�t 13ppw@"S�z�sq ~��~V�q ~ q ~�t 130ppw@$      sq ~���ʞ�q ~ q ~�t 1300ppw@$      sq ~���ʢ�q ~ q ~�t 1301ppw@$      sq ~���ʦuq ~ q ~�t 1302ppw@$      sq ~���ʪ6q ~ q ~�t 1303ppw@$      sq ~���ʭ�q ~ q ~�t 1304ppw@$      sq ~���ʱ�q ~ q ~�t 1305ppw@$      sq ~���ʵyq ~ q ~�t 1306ppw@$      sq ~���ʹ:q ~ q ~�t 1307ppw@$      sq ~���ʼ�q ~ q ~�t 1308ppw@$      sq ~������q ~ q ~�t 1309ppw@$      sq ~��~Z`q ~ q ~�t 131ppw@$      sq ~����Rq ~ q ~�t 1310ppw@$      sq ~����q ~ q ~�t 1311ppw@$      sq ~�����q ~ q ~�t 1312ppw@$      sq ~�����q ~ q ~�t 1313ppw@$      sq ~����"Vq ~ q ~�t 1314ppw@$      sq ~����&q ~ q ~�t 1315ppw@$      sq ~����)�q ~ q ~�t 1316ppw@$      sq ~����-�q ~ q ~�t 1317ppw@$      sq ~����1Zq ~ q ~�t 1318ppw@$      sq ~����5q ~ q ~�t 1319ppw@$      sq ~��~^!q ~ q ~�t 132ppw@$      sq ~���ˇ�q ~ q ~�t 1320ppw@$      sq ~���ˋrq ~ q ~�t 1321ppw@$      sq ~���ˏ3q ~ q ~�t 1322ppw@$      sq ~���˒�q ~ q ~�t 1323ppw@$      sq ~���˖�q ~ q ~�t 1324ppw@$      sq ~���˚vq ~ q ~�t 1325ppw@$      sq ~���˞7q ~ q ~�t 1326ppw@$      sq ~���ˡ�q ~ q ~�t 1327ppw@$      sq ~���˥�q ~ q ~�t 1328ppw@$      sq ~���˩zq ~ q ~�t 1329ppw@$      sq ~��~a�q ~ q ~�t 133ppw@$      sq ~�����q ~ q ~�t 1330ppw@$      sq ~������q ~ q ~�t 1331ppw@$      sq ~�����q ~ q ~�t 1332ppw@$      sq ~����Sq ~ q ~�t 1333ppw@$      sq ~����q ~ q ~�t 1334ppw@(E#�� �sq ~�����q ~ q ~�t 1335ppw@$      sq ~�����q ~ q ~�t 1336ppw@$      sq ~����Wq ~ q ~�t 1337ppw@$      sq ~����q ~ q ~�t 1338ppw@$      sq ~�����q ~ q ~�t 1339ppw@$      sq ~��~e�q ~ q ~�t 134ppw@$      sq ~����poq ~ q ~�t 1340ppw@$      sq ~����t0q ~ q ~�t 1341ppw@%����i%sq ~����w�q ~ q ~�t 1342ppw@$      sq ~����{�q ~ q ~�t 1343ppw@$      sq ~����sq ~ q ~�t 1344ppw@$      sq ~���̃4q ~ q ~�t 1345ppw@$      sq ~���̆�q ~ q ~�t 1346ppw@$      sq ~���̊�q ~ q ~�t 1347ppw@$      sq ~���̎wq ~ q ~�t 1348ppw@$      sq ~���̒8q ~ q ~�t 1349ppw@$      sq ~��~idq ~ q ~�t 135ppw@$      sq ~������q ~ q ~�t 1350ppw@$      sq ~�����q ~ q ~�t 1351ppw@$      sq ~�����Pq ~ q ~�t 1352ppw@$      sq ~�����q ~ q ~�t 1353ppw@$      sq ~������q ~ q ~�t 1354ppw@$      sq ~������q ~ q ~�t 1355ppw@$      sq ~�����Tq ~ q ~�t 1356ppw@$      sq ~�����q ~ q ~�t 1357ppw@$      sq ~�����q ~ q ~�t 1358ppw@$      sq ~�����q ~ q ~�t 1359ppw@$      sq ~��~m%q ~ q ~�t 136ppw@$      sq ~����Y-q ~ q ~�t 1360ppw@$      sq ~����\�q ~ q ~�t 1361ppw@$      sq ~����`�q ~ q ~�t 1362ppw@$      sq ~����dpq ~ q ~�t 1363ppw@$      sq ~����h1q ~ q ~�t 1364ppw@$      sq ~����k�q ~ q ~�t 1365ppw@$      sq ~����o�q ~ q ~�t 1366ppw@%���L_sq ~����stq ~ q ~�t 1367ppw@$      sq ~����w5q ~ q ~�t 1368ppw@$      sq ~����z�q ~ q ~�t 1369ppw@$      sq ~��~p�q ~ q ~�t 137ppw@$      sq ~����͌q ~ q ~�t 1370ppw@$      sq ~�����Mq ~ q ~�t 1371ppw@$      sq ~�����q ~ q ~�t 1372ppw@$      sq ~������q ~ q ~�t 1373ppw@$      sq ~����ܐq ~ q ~�t 1374ppw@$      sq ~�����Qq ~ q ~�t 1375ppw@$      sq ~�����q ~ q ~�t 1376ppw@$      sq ~������q ~ q ~�t 1377ppw@$      sq ~�����q ~ q ~�t 1378ppw@$      sq ~�����Uq ~ q ~�t 1379ppw@$      sq ~��~t�q ~ q ~�t 138ppw@$      sq ~����A�q ~ q ~�t 1380ppw@$      sq ~����E�q ~ q ~�t 1381ppw@$      sq ~����Imq ~ q ~�t 1382ppw@$      sq ~����M.q ~ q ~�t 1383ppw@$      sq ~����P�q ~ q ~�t 1384ppw@$      sq ~����T�q ~ q ~�t 1385ppw@$      sq ~����Xqq ~ q ~�t 1386ppw@$      sq ~����\2q ~ q ~�t 1387ppw@$      sq ~����_�q ~ q ~�t 1388ppw@$      sq ~����c�q ~ q ~�t 1389ppw@$      sq ~��~xhq ~ q ~�t 139ppw@$      sq ~���ζJq ~ q ~�t 1390ppw@$      sq ~���κq ~ q ~�t 1391ppw@$      sq ~���ν�q ~ q ~�t 1392ppw@$      sq ~������q ~ q ~�t 1393ppw@$      sq ~�����Nq ~ q ~�t 1394ppw@$      sq ~�����q ~ q ~�t 1395ppw@$      sq ~������q ~ q ~�t 1396ppw@$      sq ~����Бq ~ q ~�t 1397ppw@$      sq ~�����Rq ~ q ~�t 1398ppw@$      sq ~�����q ~ q ~�t 1399ppw@%�����sq ~��{^�4q ~ q ~�t 14ppw@$      sq ~��~��q ~ q ~�t 140ppw@$      sq ~���ضtq ~ q ~�t 1400ppw@$      sq ~���غ5q ~ q ~�t 1401ppw@$      sq ~���ؽ�q ~ q ~�t 1402ppw@$      sq ~������q ~ q ~�t 1403ppw@$      sq ~�����xq ~ q ~�t 1404ppw@$      sq ~�����9q ~ q ~�t 1405ppw@$      sq ~������q ~ q ~�t 1406ppw@$      sq ~����лq ~ q ~�t 1407ppw@$      sq ~�����|q ~ q ~�t 1408ppw@$      sq ~�����=q ~ q ~�t 1409ppw@$      sq ~��~οq ~ q ~�t 141ppw@$      sq ~����*�q ~ q ~�t 1410ppw@$      sq ~����.�q ~ q ~�t 1411ppw@%�ճ���sq ~����2Uq ~ q ~�t 1412ppw@$      sq ~����6q ~ q ~�t 1413ppw@$      sq ~����9�q ~ q ~�t 1414ppw@$      sq ~����=�q ~ q ~�t 1415ppw@$      sq ~����AYq ~ q ~�t 1416ppw@$      sq ~����Eq ~ q ~�t 1417ppw@$      sq ~����H�q ~ q ~�t 1418ppw@$      sq ~����L�q ~ q ~�t 1419ppw@$      sq ~��~Ҁq ~ q ~�t 142ppw@$      sq ~���ٟ2q ~ q ~�t 1420ppw@$      sq ~���٢�q ~ q ~�t 1421ppw@$      sq ~���٦�q ~ q ~�t 1422ppw@$      sq ~���٪uq ~ q ~�t 1423ppw@$      sq ~���ٮ6q ~ q ~�t 1424ppw@$      sq ~���ٱ�q ~ q ~�t 1425ppw@$      sq ~���ٵ�q ~ q ~�t 1426ppw@$      sq ~���ٹyq ~ q ~�t 1427ppw@$      sq ~���ٽ:q ~ q ~�t 1428ppw@$      sq ~������q ~ q ~�t 1429ppw@$      sq ~��~�Aq ~ q ~�t 143ppw@$      sq ~�����q ~ q ~�t 1430ppw@$      sq ~����Rq ~ q ~�t 1431ppw@$      sq ~����q ~ q ~�t 1432ppw@$      sq ~�����q ~ q ~�t 1433ppw@$      sq ~����"�q ~ q ~�t 1434ppw@$      sq ~����&Vq ~ q ~�t 1435ppw@$      sq ~����*q ~ q ~�t 1436ppw@$      sq ~����-�q ~ q ~�t 1437ppw@$      sq ~����1�q ~ q ~�t 1438ppw@$      sq ~����5Zq ~ q ~�t 1439ppw@$      sq ~��~�q ~ q ~�t 144ppw@$      sq ~���ڇ�q ~ q ~�t 1440ppw@$      sq ~���ڋ�q ~ q ~�t 1441ppw@$      sq ~���ڏrq ~ q ~�t 1442ppw@$      sq ~���ړ3q ~ q ~�t 1443ppw@$      sq ~���ږ�q ~ q ~�t 1444ppw@$      sq ~���ښ�q ~ q ~�t 1445ppw@$      sq ~���ڞvq ~ q ~�t 1446ppw@$>g�	��sq ~���ڢ7q ~ q ~�t 1447ppw@$      sq ~���ڥ�q ~ q ~�t 1448ppw@$      sq ~���ک�q ~ q ~�t 1449ppw@$      sq ~��~��q ~ q ~�t 145ppw@$      sq ~�����Oq ~ q ~�t 1450ppw@$      sq ~���� q ~ q ~�t 1451ppw@$      sq ~�����q ~ q ~�t 1452ppw@$      sq ~�����q ~ q ~�t 1453ppw@$      sq ~����Sq ~ q ~�t 1454ppw@$      sq ~����q ~ q ~�t 1455ppw@$      sq ~�����q ~ q ~�t 1456ppw@$      sq ~�����q ~ q ~�t 1457ppw@$      sq ~����Wq ~ q ~�t 1458ppw@$      sq ~����q ~ q ~�t 1459ppw@$      sq ~��~�q ~ q ~�t 146ppw@$      sq ~����p�q ~ q ~�t 1460ppw@$      sq ~����toq ~ q ~�t 1461ppw@$      sq ~����x0q ~ q ~�t 1462ppw@$      sq ~����{�q ~ q ~�t 1463ppw@$      sq ~�����q ~ q ~�t 1464ppw@$      sq ~���ۃsq ~ q ~�t 1465ppw@$      sq ~���ۇ4q ~ q ~�t 1466ppw@$      sq ~���ۊ�q ~ q ~�t 1467ppw@&      sq ~���ێ�q ~ q ~�t 1468ppw@$      sq ~���ےwq ~ q ~�t 1469ppw@$      sq ~��~�Eq ~ q ~�t 147ppw@$      sq ~�����q ~ q ~�t 1470ppw@$      sq ~������q ~ q ~�t 1471ppw@$      sq ~�����q ~ q ~�t 1472ppw@$      sq ~�����Pq ~ q ~�t 1473ppw@$      sq ~�����q ~ q ~�t 1474ppw@$      sq ~������q ~ q ~�t 1475ppw@$      sq ~������q ~ q ~�t 1476ppw@$      sq ~�����Tq ~ q ~�t 1477ppw@$      sq ~����q ~ q ~�t 1478ppw@$      sq ~�����q ~ q ~�t 1479ppw@$      sq ~��~�q ~ q ~�t 148ppw@$      sq ~����Ylq ~ q ~�t 1480ppw@$      sq ~����]-q ~ q ~�t 1481ppw@$      sq ~����`�q ~ q ~�t 1482ppw@$      sq ~����d�q ~ q ~�t 1483ppw@$      sq ~����hpq ~ q ~�t 1484ppw@$      sq ~����l1q ~ q ~�t 1485ppw@$      sq ~����o�q ~ q ~�t 1486ppw@$      sq ~����s�q ~ q ~�t 1487ppw@$      sq ~����wtq ~ q ~�t 1488ppw@$      sq ~����{5q ~ q ~�t 1489ppw@$      sq ~��~��q ~ q ~�t 149ppw@'��D�;^sq ~������q ~ q ~�t 1490ppw@$      sq ~����ьq ~ q ~�t 1491ppw@$      sq ~�����Mq ~ q ~�t 1492ppw@$      sq ~�����q ~ q ~�t 1493ppw@$      sq ~������q ~ q ~�t 1494ppw@$      sq ~������q ~ q ~�t 1495ppw@$      sq ~�����Qq ~ q ~�t 1496ppw@#�k�(&sq ~�����q ~ q ~�t 1497ppw@$      sq ~������q ~ q ~�t 1498ppw@$      sq ~�����q ~ q ~�t 1499ppw@$      sq ~��{_ �q ~ q ~�t 15ppw@@��Ъ�sq ~��~?]q ~ q ~�t 150ppw@$      sq ~������q ~ q ~�t 1500ppw@$      sq ~����Ѷq ~ q ~�t 1501ppw@$      sq ~�����wq ~ q ~�t 1502ppw@$      sq ~�����8q ~ q ~�t 1503ppw@$      sq ~������q ~ q ~�t 1504ppw@$      sq ~�����q ~ q ~�t 1505ppw@$      sq ~�����{q ~ q ~�t 1506ppw@$      sq ~�����<q ~ q ~�t 1507ppw@$      sq ~������q ~ q ~�t 1508ppw@$      sq ~�����q ~ q ~�t 1509ppw@$      sq ~��~Cq ~ q ~�t 151ppw@$      sq ~����BTq ~ q ~�t 1510ppw@$      sq ~����Fq ~ q ~�t 1511ppw@$      sq ~����I�q ~ q ~�t 1512ppw@$      sq ~����M�q ~ q ~�t 1513ppw@$      sq ~����QXq ~ q ~�t 1514ppw@$      sq ~����Uq ~ q ~�t 1515ppw@$      sq ~����X�q ~ q ~�t 1516ppw@$      sq ~����\�q ~ q ~�t 1517ppw@$      sq ~����`\q ~ q ~�t 1518ppw@$      sq ~����dq ~ q ~�t 1519ppw@$      sq ~��~F�q ~ q ~�t 152ppw@$      sq ~���綳q ~ q ~�t 1520ppw@$      sq ~����tq ~ q ~�t 1521ppw@$      sq ~����5q ~ q ~�t 1522ppw@$      sq ~������q ~ q ~�t 1523ppw@$      sq ~����ŷq ~ q ~�t 1524ppw@$      sq ~�����xq ~ q ~�t 1525ppw@$      sq ~�����9q ~ q ~�t 1526ppw@$      sq ~������q ~ q ~�t 1527ppw@$      sq ~����Իq ~ q ~�t 1528ppw@$      sq ~�����|q ~ q ~�t 1529ppw@$      sq ~��~J�q ~ q ~�t 153ppw@$      sq ~����+q ~ q ~�t 1530ppw@$      sq ~����.�q ~ q ~�t 1531ppw@$      sq ~����2�q ~ q ~�t 1532ppw@$      sq ~����6Uq ~ q ~�t 1533ppw@$      sq ~����:q ~ q ~�t 1534ppw@$      sq ~����=�q ~ q ~�t 1535ppw@$      sq ~����A�q ~ q ~�t 1536ppw@$      sq ~����EYq ~ q ~�t 1537ppw@$      sq ~����Iq ~ q ~�t 1538ppw@$      sq ~����L�q ~ q ~�t 1539ppw@$      sq ~��~Naq ~ q ~�t 154ppw@$      sq ~����qq ~ q ~�t 1540ppw@$      sq ~����2q ~ q ~�t 1541ppw@$      sq ~�����q ~ q ~�t 1542ppw@$      sq ~���誴q ~ q ~�t 1543ppw@$      sq ~����uq ~ q ~�t 1544ppw@$      sq ~����6q ~ q ~�t 1545ppw@$      sq ~�����q ~ q ~�t 1546ppw@$      sq ~���蹸q ~ q ~�t 1547ppw@%�)hGtsq ~����yq ~ q ~�t 1548ppw@$      sq ~�����:q ~ q ~�t 1549ppw@$      sq ~��~R"q ~ q ~�t 155ppw@$      sq ~�����q ~ q ~�t 1550ppw@$      sq ~�����q ~ q ~�t 1551ppw@$      sq ~����Rq ~ q ~�t 1552ppw@$      sq ~����q ~ q ~�t 1553ppw@$      sq ~����"�q ~ q ~�t 1554ppw@$      sq ~����&�q ~ q ~�t 1555ppw@$      sq ~����*Vq ~ q ~�t 1556ppw@$      sq ~����.q ~ q ~�t 1557ppw@$      sq ~����1�q ~ q ~�t 1558ppw@$      sq ~����5�q ~ q ~�t 1559ppw@$      sq ~��~U�q ~ q ~�t 156ppw@$      sq ~����/q ~ q ~�t 1560ppw@$      sq ~�����q ~ q ~�t 1561ppw@$      sq ~���鏱q ~ q ~�t 1562ppw@$      sq ~����rq ~ q ~�t 1563ppw@$      sq ~����3q ~ q ~�t 1564ppw@$      sq ~�����q ~ q ~�t 1565ppw@$      sq ~���鞵q ~ q ~�t 1566ppw@$      sq ~����vq ~ q ~�t 1567ppw@$      sq ~����7q ~ q ~�t 1568ppw@$      sq ~�����q ~ q ~�t 1569ppw@$      sq ~��~Y�q ~ q ~�t 157ppw@$      sq ~������q ~ q ~�t 1570ppw@$      sq ~���� Oq ~ q ~�t 1571ppw@$      sq ~����q ~ q ~�t 1572ppw@$      sq ~�����q ~ q ~�t 1573ppw@$      sq ~�����q ~ q ~�t 1574ppw@$      sq ~����Sq ~ q ~�t 1575ppw@$      sq ~����q ~ q ~�t 1576ppw@$      sq ~�����q ~ q ~�t 1577ppw@$      sq ~�����q ~ q ~�t 1578ppw@$      sq ~����Wq ~ q ~�t 1579ppw@$      sq ~��~]eq ~ q ~�t 158ppw@$      sq ~����p�q ~ q ~�t 1580ppw@$      sq ~����t�q ~ q ~�t 1581ppw@$      sq ~����xoq ~ q ~�t 1582ppw@$      sq ~����|0q ~ q ~�t 1583ppw@$      sq ~�����q ~ q ~�t 1584ppw@$      sq ~���ꃲq ~ q ~�t 1585ppw@$      sq ~����sq ~ q ~�t 1586ppw@$      sq ~����4q ~ q ~�t 1587ppw@$      sq ~�����q ~ q ~�t 1588ppw@$      sq ~���꒶q ~ q ~�t 1589ppw@$      sq ~��~a&q ~ q ~�t 159ppw@$      sq ~�����Lq ~ q ~�t 1590ppw@$      sq ~�����q ~ q ~�t 1591ppw@$      sq ~������q ~ q ~�t 1592ppw@$      sq ~������q ~ q ~�t 1593ppw@$      sq ~�����Pq ~ q ~�t 1594ppw@$      sq ~�����q ~ q ~�t 1595ppw@$      sq ~������q ~ q ~�t 1596ppw@$      sq ~������q ~ q ~�t 1597ppw@$      sq ~����Tq ~ q ~�t 1598ppw@$      sq ~����q ~ q ~�t 1599ppw@$      sq ~��{_�q ~ q ~�t 16ppw@$      sq ~��~��q ~ q ~�t 160ppw@$      sq ~�����vq ~ q ~�t 1600ppw@$      sq ~�����7q ~ q ~�t 1601ppw@$      sq ~������q ~ q ~�t 1602ppw@$      sq ~�����q ~ q ~�t 1603ppw@$      sq ~�����zq ~ q ~�t 1604ppw@$      sq ~�����;q ~ q ~�t 1605ppw@$      sq ~������q ~ q ~�t 1606ppw@$      sq ~������q ~ q ~�t 1607ppw@$      sq ~����~q ~ q ~�t 1608ppw@$      sq ~����?q ~ q ~�t 1609ppw@$      sq ~��~�}q ~ q ~�t 161ppw@$      sq ~����Y�q ~ q ~�t 1610ppw@$      sq ~����]�q ~ q ~�t 1611ppw@$      sq ~����aWq ~ q ~�t 1612ppw@$      sq ~����eq ~ q ~�t 1613ppw@$      sq ~����h�q ~ q ~�t 1614ppw@$      sq ~����l�q ~ q ~�t 1615ppw@$      sq ~����p[q ~ q ~�t 1616ppw@$      sq ~����tq ~ q ~�t 1617ppw@$      sq ~����w�q ~ q ~�t 1618ppw@$      sq ~����{�q ~ q ~�t 1619ppw@$      sq ~��~�>q ~ q ~�t 162ppw@$      sq ~�����4q ~ q ~�t 1620ppw@$      sq ~������q ~ q ~�t 1621ppw@$      sq ~����նq ~ q ~�t 1622ppw@$      sq ~�����wq ~ q ~�t 1623ppw@$      sq ~�����8q ~ q ~�t 1624ppw@$      sq ~������q ~ q ~�t 1625ppw@$      sq ~�����q ~ q ~�t 1626ppw@$      sq ~�����{q ~ q ~�t 1627ppw@$      sq ~�����<q ~ q ~�t 1628ppw@$      sq ~������q ~ q ~�t 1629ppw@$      sq ~��~��q ~ q ~�t 163ppw@$      sq ~����B�q ~ q ~�t 1630ppw@$      sq ~����FTq ~ q ~�t 1631ppw@$      sq ~����Jq ~ q ~�t 1632ppw@$      sq ~����M�q ~ q ~�t 1633ppw@$      sq ~����Q�q ~ q ~�t 1634ppw@$      sq ~����UXq ~ q ~�t 1635ppw@$      sq ~����Yq ~ q ~�t 1636ppw@$      sq ~����\�q ~ q ~�t 1637ppw@$      sq ~����`�q ~ q ~�t 1638ppw@$      sq ~����d\q ~ q ~�t 1639ppw@$      sq ~��~��q ~ q ~�t 164ppw@$      sq ~������q ~ q ~�t 1640ppw@$      sq ~������q ~ q ~�t 1641ppw@$      sq ~�����tq ~ q ~�t 1642ppw@$      sq ~�����5q ~ q ~�t 1643ppw@$      sq ~������q ~ q ~�t 1644ppw@$      sq ~����ɷq ~ q ~�t 1645ppw@$      sq ~�����xq ~ q ~�t 1646ppw@$      sq ~�����9q ~ q ~�t 1647ppw@$      sq ~������q ~ q ~�t 1648ppw@$      sq ~����ػq ~ q ~�t 1649ppw@$      sq ~��~Ɓq ~ q ~�t 165ppw@$      sq ~����+Qq ~ q ~�t 1650ppw@$      sq ~����/q ~ q ~�t 1651ppw@$      sq ~����2�q ~ q ~�t 1652ppw@$      sq ~����6�q ~ q ~�t 1653ppw@$      sq ~����:Uq ~ q ~�t 1654ppw@$      sq ~����>q ~ q ~�t 1655ppw@$      sq ~����A�q ~ q ~�t 1656ppw@$      sq ~����E�q ~ q ~�t 1657ppw@$      sq ~����IYq ~ q ~�t 1658ppw@$      sq ~����Mq ~ q ~�t 1659ppw@$      sq ~��~�Bq ~ q ~�t 166ppw@$      sq ~������q ~ q ~�t 1660ppw@$      sq ~�����qq ~ q ~�t 1661ppw@$      sq ~�����2q ~ q ~�t 1662ppw@$      sq ~������q ~ q ~�t 1663ppw@$      sq ~������q ~ q ~�t 1664ppw@&5�k�sq ~�����uq ~ q ~�t 1665ppw@$      sq ~�����6q ~ q ~�t 1666ppw@$      sq ~������q ~ q ~�t 1667ppw@$      sq ~������q ~ q ~�t 1668ppw@$      sq ~�����yq ~ q ~�t 1669ppw@$      sq ~��~�q ~ q ~�t 167ppw@$      sq ~����q ~ q ~�t 1670ppw@$      sq ~�����q ~ q ~�t 1671ppw@$      sq ~�����q ~ q ~�t 1672ppw@$      sq ~����Rq ~ q ~�t 1673ppw@$      sq ~����#q ~ q ~�t 1674ppw@$      sq ~����&�q ~ q ~�t 1675ppw@$      sq ~����*�q ~ q ~�t 1676ppw@$      sq ~����.Vq ~ q ~�t 1677ppw@$      sq ~����2q ~ q ~�t 1678ppw@$      sq ~����5�q ~ q ~�t 1679ppw@$      sq ~��~��q ~ q ~�t 168ppw@$      sq ~�����nq ~ q ~�t 1680ppw@$      sq ~�����/q ~ q ~�t 1681ppw@$      sq ~������q ~ q ~�t 1682ppw@$      sq ~������q ~ q ~�t 1683ppw@$      sq ~�����rq ~ q ~�t 1684ppw@$      sq ~�����3q ~ q ~�t 1685ppw@$      sq ~������q ~ q ~�t 1686ppw@$      sq ~������q ~ q ~�t 1687ppw@$O,5/*�sq ~�����vq ~ q ~�t 1688ppw@$      sq ~�����7q ~ q ~�t 1689ppw@$      sq ~��~Յq ~ q ~�t 169ppw@$      sq ~������q ~ q ~�t 1690ppw@$      sq ~���� �q ~ q ~�t 1691ppw@$      sq ~����Oq ~ q ~�t 1692ppw@$      sq ~����q ~ q ~�t 1693ppw@$      sq ~�����q ~ q ~�t 1694ppw@$      sq ~�����q ~ q ~�t 1695ppw@$      sq ~����Sq ~ q ~�t 1696ppw@$      sq ~����q ~ q ~�t 1697ppw@$      sq ~�����q ~ q ~�t 1698ppw@$      sq ~�����q ~ q ~�t 1699ppw@$      sq ~��{_wq ~ q ~�t 17ppw@/��m�6 sq ~��~(q ~ q ~�t 170ppw@$      sq ~�����q ~ q ~�t 1700ppw@$      sq ~��� �q ~ q ~�t 1701ppw@$      sq ~���yq ~ q ~�t 1702ppw@$      sq ~���:q ~ q ~�t 1703ppw@$      sq ~����q ~ q ~�t 1704ppw@$      sq ~����q ~ q ~�t 1705ppw@$      sq ~���}q ~ q ~�t 1706ppw@$      sq ~���>q ~ q ~�t 1707ppw@$      sq ~����q ~ q ~�t 1708ppw@$      sq ~����q ~ q ~�t 1709ppw@$      sq ~��~+�q ~ q ~�t 171ppw@$      sq ~���qVq ~ q ~�t 1710ppw@$      sq ~���uq ~ q ~�t 1711ppw@$      sq ~���x�q ~ q ~�t 1712ppw@$      sq ~���|�q ~ q ~�t 1713ppw@$      sq ~����Zq ~ q ~�t 1714ppw@$      sq ~����q ~ q ~�t 1715ppw@$      sq ~�����q ~ q ~�t 1716ppw@$      sq ~�����q ~ q ~�t 1717ppw@$      sq ~����^q ~ q ~�t 1718ppw@$      sq ~����q ~ q ~�t 1719ppw@$      sq ~��~/�q ~ q ~�t 172ppw@$      sq ~����q ~ q ~�t 1720ppw@$      sq ~����vq ~ q ~�t 1721ppw@$      sq ~����7q ~ q ~�t 1722ppw@$      sq ~�����q ~ q ~�t 1723ppw@$      sq ~�����q ~ q ~�t 1724ppw@$      sq ~����zq ~ q ~�t 1725ppw@"D�^���sq ~����;q ~ q ~�t 1726ppw@$      sq ~�����q ~ q ~�t 1727ppw@$      sq ~����q ~ q ~�t 1728ppw@$      sq ~���~q ~ q ~�t 1729ppw@$      sq ~��~3^q ~ q ~�t 173ppw@$      sq ~���Zq ~ q ~�t 1730ppw@$      sq ~���]�q ~ q ~�t 1731ppw@$      sq ~���a�q ~ q ~�t 1732ppw@$      sq ~���eWq ~ q ~�t 1733ppw@$      sq ~���iq ~ q ~�t 1734ppw@$      sq ~���l�q ~ q ~�t 1735ppw@$      sq ~���p�q ~ q ~�t 1736ppw@$      sq ~���t[q ~ q ~�t 1737ppw@$      sq ~���xq ~ q ~�t 1738ppw@$      sq ~���{�q ~ q ~�t 1739ppw@$      sq ~��~7q ~ q ~�t 174ppw@$      sq ~����sq ~ q ~�t 1740ppw@$      sq ~����4q ~ q ~�t 1741ppw@$      sq ~�����q ~ q ~�t 1742ppw@$      sq ~���ٶq ~ q ~�t 1743ppw@$      sq ~����wq ~ q ~�t 1744ppw@$      sq ~����8q ~ q ~�t 1745ppw@$��&�sq ~�����q ~ q ~�t 1746ppw@$      sq ~����q ~ q ~�t 1747ppw@$      sq ~����{q ~ q ~�t 1748ppw@$      sq ~����<q ~ q ~�t 1749ppw@$      sq ~��~:�q ~ q ~�t 175ppw@$      sq ~���B�q ~ q ~�t 1750ppw@$      sq ~���F�q ~ q ~�t 1751ppw@$      sq ~���JTq ~ q ~�t 1752ppw@$      sq ~���Nq ~ q ~�t 1753ppw@$      sq ~���Q�q ~ q ~�t 1754ppw@$      sq ~���U�q ~ q ~�t 1755ppw@$      sq ~���YXq ~ q ~�t 1756ppw@$      sq ~���]q ~ q ~�t 1757ppw@$      sq ~���`�q ~ q ~�t 1758ppw@$      sq ~���d�q ~ q ~�t 1759ppw@$      sq ~��~>�q ~ q ~�t 176ppw@$      sq ~����1q ~ q ~�t 1760ppw@$      sq ~�����q ~ q ~�t 1761ppw@$      sq ~�����q ~ q ~�t 1762ppw@$      sq ~����tq ~ q ~�t 1763ppw@$      sq ~����5q ~ q ~�t 1764ppw@$      sq ~�����q ~ q ~�t 1765ppw@$      sq ~���ͷq ~ q ~�t 1766ppw@$      sq ~����xq ~ q ~�t 1767ppw@$      sq ~����9q ~ q ~�t 1768ppw@$      sq ~�����q ~ q ~�t 1769ppw@$      sq ~��~Bbq ~ q ~�t 177ppw@$      sq ~���+�q ~ q ~�t 1770ppw@$      sq ~���/Qq ~ q ~�t 1771ppw@$      sq ~���3q ~ q ~�t 1772ppw@$      sq ~���6�q ~ q ~�t 1773ppw@$      sq ~���:�q ~ q ~�t 1774ppw@$      sq ~���>Uq ~ q ~�t 1775ppw@$      sq ~���Bq ~ q ~�t 1776ppw@$      sq ~���E�q ~ q ~�t 1777ppw@$      sq ~���I�q ~ q ~�t 1778ppw@ � ��'�sq ~���MYq ~ q ~�t 1779ppw@$      sq ~��~F#q ~ q ~�t 178ppw@$      sq ~�����q ~ q ~�t 1780ppw@$      sq ~�����q ~ q ~�t 1781ppw@$      sq ~����qq ~ q ~�t 1782ppw@$      sq ~����2q ~ q ~�t 1783ppw@$      sq ~�����q ~ q ~�t 1784ppw@$      sq ~�����q ~ q ~�t 1785ppw@$      sq ~����uq ~ q ~�t 1786ppw@$      sq ~����6q ~ q ~�t 1787ppw@$      sq ~�����q ~ q ~�t 1788ppw@$      sq ~�����q ~ q ~�t 1789ppw@#y�Ƚsq ~��~I�q ~ q ~�t 179ppw@$      sq ~���Nq ~ q ~�t 1790ppw@$      sq ~���q ~ q ~�t 1791ppw@$      sq ~����q ~ q ~�t 1792ppw@$      sq ~����q ~ q ~�t 1793ppw@$      sq ~���#Rq ~ q ~�t 1794ppw@$      sq ~���'q ~ q ~�t 1795ppw@$      sq ~���*�q ~ q ~�t 1796ppw@$      sq ~���.�q ~ q ~�t 1797ppw@33���H?sq ~���2Vq ~ q ~�t 1798ppw@$      sq ~���6q ~ q ~�t 1799ppw@$      sq ~��{_8q ~ q ~�t 18ppw@ 5�v� |sq ~��~�zq ~ q ~�t 180ppw@$      sq ~���xq ~ q ~�t 1800ppw@$      sq ~���9q ~ q ~�t 1801ppw@$      sq ~����q ~ q ~�t 1802ppw@$      sq ~����q ~ q ~�t 1803ppw@$      sq ~���#|q ~ q ~�t 1804ppw@$      sq ~���'=q ~ q ~�t 1805ppw@$      sq ~���*�q ~ q ~�t 1806ppw@$      sq ~���.�q ~ q ~�t 1807ppw@$      sq ~���2�q ~ q ~�t 1808ppw@$      sq ~���6Aq ~ q ~�t 1809ppw@$      sq ~��~�;q ~ q ~�t 181ppw@$      sq ~�����q ~ q ~�t 1810ppw@$      sq ~�����q ~ q ~�t 1811ppw@$      sq ~����Yq ~ q ~�t 1812ppw@%�]�7�sq ~����q ~ q ~�t 1813ppw@$      sq ~�����q ~ q ~�t 1814ppw@$      sq ~�����q ~ q ~�t 1815ppw@$      sq ~����]q ~ q ~�t 1816ppw@#�)6I�sq ~����q ~ q ~�t 1817ppw@$      sq ~�����q ~ q ~�t 1818ppw@$      sq ~�����q ~ q ~�t 1819ppw@$      sq ~��~��q ~ q ~�t 182ppw@$      sq ~����6q ~ q ~�t 1820ppw@$      sq ~��� �q ~ q ~�t 1821ppw@$      sq ~����q ~ q ~�t 1822ppw@$      sq ~���yq ~ q ~�t 1823ppw@$      sq ~���:q ~ q ~�t 1824ppw@$      sq ~����q ~ q ~�t 1825ppw@$      sq ~����q ~ q ~�t 1826ppw@$      sq ~���}q ~ q ~�t 1827ppw@$      sq ~���>q ~ q ~�t 1828ppw@$      sq ~����q ~ q ~�t 1829ppw@%�ذ�|
sq ~��~��q ~ q ~�t 183ppw@$      sq ~���q�q ~ q ~�t 1830ppw@$      sq ~���uVq ~ q ~�t 1831ppw@$      sq ~���yq ~ q ~�t 1832ppw@$      sq ~���|�q ~ q ~�t 1833ppw@$      sq ~�����q ~ q ~�t 1834ppw@$      sq ~����Zq ~ q ~�t 1835ppw@$      sq ~����q ~ q ~�t 1836ppw@$      sq ~�����q ~ q ~�t 1837ppw@$      sq ~�����q ~ q ~�t 1838ppw@$      sq ~����^q ~ q ~�t 1839ppw@$      sq ~��~�~q ~ q ~�t 184ppw@$      sq ~�����q ~ q ~�t 1840ppw@$      sq ~����q ~ q ~�t 1841ppw@$      sq ~����vq ~ q ~�t 1842ppw@$      sq ~����7q ~ q ~�t 1843ppw@$      sq ~�����q ~ q ~�t 1844ppw@$      sq ~�����q ~ q ~�t 1845ppw@$      sq ~����zq ~ q ~�t 1846ppw@#�{�߇�sq ~��� ;q ~ q ~�t 1847ppw@$      sq ~����q ~ q ~�t 1848ppw@$      sq ~����q ~ q ~�t 1849ppw@$      sq ~��~�?q ~ q ~�t 185ppw@$      sq ~���ZSq ~ q ~�t 1850ppw@$      sq ~���^q ~ q ~�t 1851ppw@$      sq ~���a�q ~ q ~�t 1852ppw@$      sq ~���e�q ~ q ~�t 1853ppw@$      sq ~���iWq ~ q ~�t 1854ppw@$      sq ~���mq ~ q ~�t 1855ppw@$      sq ~���p�q ~ q ~�t 1856ppw@$      sq ~���t�q ~ q ~�t 1857ppw@$      sq ~���x[q ~ q ~�t 1858ppw@$      sq ~���|q ~ q ~�t 1859ppw@$      sq ~��~� q ~ q ~�t 186ppw@$      sq ~���βq ~ q ~�t 1860ppw@$      sq ~����sq ~ q ~�t 1861ppw@$      sq ~����4q ~ q ~�t 1862ppw@$      sq ~�����q ~ q ~�t 1863ppw@$      sq ~���ݶq ~ q ~�t 1864ppw@$      sq ~����wq ~ q ~�t 1865ppw@$      sq ~����8q ~ q ~�t 1866ppw@$      sq ~�����q ~ q ~�t 1867ppw@$      sq ~����q ~ q ~�t 1868ppw@$      sq ~����{q ~ q ~�t 1869ppw@$      sq ~��~��q ~ q ~�t 187ppw@$      sq ~���Cq ~ q ~�t 1870ppw@$      sq ~���F�q ~ q ~�t 1871ppw@$      sq ~���J�q ~ q ~�t 1872ppw@$      sq ~���NTq ~ q ~�t 1873ppw@$      sq ~���Rq ~ q ~�t 1874ppw@$      sq ~���U�q ~ q ~�t 1875ppw@$      sq ~���Y�q ~ q ~�t 1876ppw@$      sq ~���]Xq ~ q ~�t 1877ppw@$      sq ~���aq ~ q ~�t 1878ppw@$      sq ~���d�q ~ q ~�t 1879ppw@"D�^�v.sq ~��~��q ~ q ~�t 188ppw@$      sq ~����pq ~ q ~�t 1880ppw@$      sq ~����1q ~ q ~�t 1881ppw@$      sq ~�����q ~ q ~�t 1882ppw@$      sq ~���³q ~ q ~�t 1883ppw@$      sq ~����tq ~ q ~�t 1884ppw@$)�xjysq ~����5q ~ q ~�t 1885ppw@$      sq ~�����q ~ q ~�t 1886ppw@$      sq ~���ѷq ~ q ~�t 1887ppw@$      sq ~����xq ~ q ~�t 1888ppw@$      sq ~����9q ~ q ~�t 1889ppw@$      sq ~��~�Cq ~ q ~�t 189ppw@$      sq ~���+�q ~ q ~�t 1890ppw@$      sq ~���/�q ~ q ~�t 1891ppw@$      sq ~���3Qq ~ q ~�t 1892ppw@$      sq ~���7q ~ q ~�t 1893ppw@$      sq ~���:�q ~ q ~�t 1894ppw@$      sq ~���>�q ~ q ~�t 1895ppw@$      sq ~���BUq ~ q ~�t 1896ppw@$      sq ~���Fq ~ q ~�t 1897ppw@$      sq ~���I�q ~ q ~�t 1898ppw@$      sq ~���M�q ~ q ~�t 1899ppw@$      sq ~��{_�q ~ q ~�t 19ppw@$      sq ~��~�q ~ q ~�t 190ppw@$      sq ~���+�q ~ q ~�t 1900ppw@$      sq ~���/�q ~ q ~�t 1901ppw@$      sq ~���3{q ~ q ~�t 1902ppw@$      sq ~���7<q ~ q ~�t 1903ppw@$      sq ~���:�q ~ q ~�t 1904ppw@$      sq ~���>�q ~ q ~�t 1905ppw@$      sq ~���Bq ~ q ~�t 1906ppw@$      sq ~���F@q ~ q ~�t 1907ppw@$      sq ~���Jq ~ q ~�t 1908ppw@$      sq ~���M�q ~ q ~�t 1909ppw@$      sq ~��~�q ~ q ~�t 191ppw@$      sq ~����Xq ~ q ~�t 1910ppw@$      sq ~����q ~ q ~�t 1911ppw@$      sq ~�����q ~ q ~�t 1912ppw@$      sq ~�����q ~ q ~�t 1913ppw@$      sq ~����\q ~ q ~�t 1914ppw@$      sq ~����q ~ q ~�t 1915ppw@$      sq ~�����q ~ q ~�t 1916ppw@$      sq ~�����q ~ q ~�t 1917ppw@$      sq ~����`q ~ q ~�t 1918ppw@$      sq ~����!q ~ q ~�t 1919ppw@$      sq ~��~[q ~ q ~�t 192ppw@$      sq ~��� �q ~ q ~�t 1920ppw@$      sq ~��� xq ~ q ~�t 1921ppw@$      sq ~��� 9q ~ q ~�t 1922ppw@$      sq ~��� �q ~ q ~�t 1923ppw@$      sq ~��� #�q ~ q ~�t 1924ppw@$      sq ~��� '|q ~ q ~�t 1925ppw@$      sq ~��� +=q ~ q ~�t 1926ppw@$      sq ~��� .�q ~ q ~�t 1927ppw@$      sq ~��� 2�q ~ q ~�t 1928ppw@$      sq ~��� 6�q ~ q ~�t 1929ppw@$      sq ~��~q ~ q ~�t 193ppw@" ��C�sq ~��� �q ~ q ~�t 1930ppw@$      sq ~��� ��q ~ q ~�t 1931ppw@$      sq ~��� ��q ~ q ~�t 1932ppw@$      sq ~��� �Yq ~ q ~�t 1933ppw@$      sq ~��� �q ~ q ~�t 1934ppw@$      sq ~��� ��q ~ q ~�t 1935ppw@$      sq ~��� ��q ~ q ~�t 1936ppw@$      sq ~��� �]q ~ q ~�t 1937ppw@#�pi[��sq ~��� �q ~ q ~�t 1938ppw@$      sq ~��� ��q ~ q ~�t 1939ppw@$      sq ~��~�q ~ q ~�t 194ppw@$      sq ~��� �uq ~ q ~�t 1940ppw@$      sq ~���!6q ~ q ~�t 1941ppw@$      sq ~���!�q ~ q ~�t 1942ppw@$      sq ~���!�q ~ q ~�t 1943ppw@$      sq ~���!yq ~ q ~�t 1944ppw@$      sq ~���!:q ~ q ~�t 1945ppw@$      sq ~���!�q ~ q ~�t 1946ppw@$      sq ~���!�q ~ q ~�t 1947ppw@$      sq ~���!}q ~ q ~�t 1948ppw@$      sq ~���!>q ~ q ~�t 1949ppw@$      sq ~��~#�q ~ q ~�t 195ppw@$      sq ~���!q�q ~ q ~�t 1950ppw@$      sq ~���!u�q ~ q ~�t 1951ppw@$      sq ~���!yVq ~ q ~�t 1952ppw@$      sq ~���!}q ~ q ~�t 1953ppw@$      sq ~���!��q ~ q ~�t 1954ppw@#��<U�+sq ~���!��q ~ q ~�t 1955ppw@$      sq ~���!�Zq ~ q ~�t 1956ppw@$      sq ~���!�q ~ q ~�t 1957ppw@$      sq ~���!��q ~ q ~�t 1958ppw@$      sq ~���!��q ~ q ~�t 1959ppw@$      sq ~��~'_q ~ q ~�t 196ppw@$      sq ~���!�3q ~ q ~�t 1960ppw@$      sq ~���!��q ~ q ~�t 1961ppw@$      sq ~���!�q ~ q ~�t 1962ppw@$      sq ~���!�vq ~ q ~�t 1963ppw@$      sq ~���!�7q ~ q ~�t 1964ppw@$      sq ~���!��q ~ q ~�t 1965ppw@$      sq ~���!��q ~ q ~�t 1966ppw@$      sq ~���" zq ~ q ~�t 1967ppw@$      sq ~���";q ~ q ~�t 1968ppw@$      sq ~���"�q ~ q ~�t 1969ppw@$      sq ~��~+ q ~ q ~�t 197ppw@$      sq ~���"Z�q ~ q ~�t 1970ppw@$      sq ~���"^Sq ~ q ~�t 1971ppw@$      sq ~���"bq ~ q ~�t 1972ppw@$      sq ~���"e�q ~ q ~�t 1973ppw@$      sq ~���"i�q ~ q ~�t 1974ppw@$      sq ~���"mWq ~ q ~�t 1975ppw@$      sq ~���"qq ~ q ~�t 1976ppw@$      sq ~���"t�q ~ q ~�t 1977ppw@$��3�sq ~���"x�q ~ q ~�t 1978ppw@$      sq ~���"|[q ~ q ~�t 1979ppw@$      sq ~��~.�q ~ q ~�t 198ppw@$      sq ~���"��q ~ q ~�t 1980ppw@$      sq ~���"Ҳq ~ q ~�t 1981ppw@$      sq ~���"�sq ~ q ~�t 1982ppw@$      sq ~���"�4q ~ q ~�t 1983ppw@$      sq ~���"��q ~ q ~�t 1984ppw@$      sq ~���"�q ~ q ~�t 1985ppw@$      sq ~���"�wq ~ q ~�t 1986ppw@$      sq ~���"�8q ~ q ~�t 1987ppw@$      sq ~���"��q ~ q ~�t 1988ppw@$      sq ~���"�q ~ q ~�t 1989ppw@$      sq ~��~2�q ~ q ~�t 199ppw@$      sq ~���#CPq ~ q ~�t 1990ppw@$      sq ~���#Gq ~ q ~�t 1991ppw@/�Z=�ݎsq ~���#J�q ~ q ~�t 1992ppw@$      sq ~���#N�q ~ q ~�t 1993ppw@$      sq ~���#RTq ~ q ~�t 1994ppw@$      sq ~���#Vq ~ q ~�t 1995ppw@$      sq ~���#Y�q ~ q ~�t 1996ppw@$      sq ~���#]�q ~ q ~�t 1997ppw@$      sq ~���#aXq ~ q ~�t 1998ppw@$      sq ~���#eq ~ q ~�t 1999ppw@$      sq ~��{H��q ~ q ~�t 2ppw@$      sq ~��{_b�q ~ q ~�t 20ppw@1t�ܑD�sq ~��~q ~ q ~�t 200ppw@$      sq ~���U1q ~ q ~�t 2000ppw@$      sq ~���U4�q ~ q ~�t 2001ppw@$      sq ~���U8�q ~ q ~�t 2002ppw@$      sq ~���U<Rq ~ q ~�t 2003ppw@$      sq ~���U@q ~ q ~�t 2004ppw@$      sq ~���UC�q ~ q ~�t 2005ppw@$      sq ~���UG�q ~ q ~�t 2006ppw@$      sq ~���UKVq ~ q ~�t 2007ppw@$      sq ~���UOq ~ q ~�t 2008ppw@$      sq ~���UR�q ~ q ~�t 2009ppw@$      sq ~��~�q ~ q ~�t 201ppw@$      sq ~���U�nq ~ q ~�t 2010ppw@$      sq ~���U�/q ~ q ~�t 2011ppw@$      sq ~���U��q ~ q ~�t 2012ppw@$      sq ~���U��q ~ q ~�t 2013ppw@$      sq ~���U�rq ~ q ~�t 2014ppw@$      sq ~���U�3q ~ q ~�t 2015ppw@$      sq ~���U��q ~ q ~�t 2016ppw@$      sq ~���U��q ~ q ~�t 2017ppw@$      sq ~���U�vq ~ q ~�t 2018ppw@$      sq ~���U�7q ~ q ~�t 2019ppw@$      sq ~��~�q ~ q ~�t 202ppw@$      sq ~���V�q ~ q ~�t 2020ppw@$      sq ~���V�q ~ q ~�t 2021ppw@$      sq ~���V!Oq ~ q ~�t 2022ppw@$      sq ~���V%q ~ q ~�t 2023ppw@$      sq ~���V(�q ~ q ~�t 2024ppw@$      sq ~���V,�q ~ q ~�t 2025ppw@$      sq ~���V0Sq ~ q ~�t 2026ppw@$      sq ~���V4q ~ q ~�t 2027ppw@$      sq ~���V7�q ~ q ~�t 2028ppw@$      sq ~���V;�q ~ q ~�t 2029ppw@$      sq ~��~Fq ~ q ~�t 203ppw@$      sq ~���V�,q ~ q ~�t 2030ppw@$      sq ~���V��q ~ q ~�t 2031ppw@$      sq ~���V��q ~ q ~�t 2032ppw@$      sq ~���V�oq ~ q ~�t 2033ppw@$      sq ~���V�0q ~ q ~�t 2034ppw@$      sq ~���V��q ~ q ~�t 2035ppw@$      sq ~���V��q ~ q ~�t 2036ppw@$      sq ~���V�sq ~ q ~�t 2037ppw@$      sq ~���V�4q ~ q ~�t 2038ppw@$      sq ~���V��q ~ q ~�t 2039ppw@$      sq ~��~ q ~ q ~�t 204ppw@$      sq ~���W�q ~ q ~�t 2040ppw@$      sq ~���WLq ~ q ~�t 2041ppw@$      sq ~���W
q ~ q ~�t 2042ppw@$      sq ~���W�q ~ q ~�t 2043ppw@$      sq ~���W�q ~ q ~�t 2044ppw@$      sq ~���WPq ~ q ~�t 2045ppw@$      sq ~���Wq ~ q ~�t 2046ppw@$      sq ~���W�q ~ q ~�t 2047ppw@$      sq ~���W �q ~ q ~�t 2048ppw@$      sq ~���W$Tq ~ q ~�t 2049ppw@$      sq ~��~#�q ~ q ~�t 205ppw@$      sq ~���Wv�q ~ q ~�t 2050ppw@$      sq ~���Wz�q ~ q ~�t 2051ppw@$      sq ~���W~lq ~ q ~�t 2052ppw@$      sq ~���W�-q ~ q ~�t 2053ppw@$      sq ~���W��q ~ q ~�t 2054ppw@$      sq ~���W��q ~ q ~�t 2055ppw@$      sq ~���W�pq ~ q ~�t 2056ppw@$      sq ~���W�1q ~ q ~�t 2057ppw@$      sq ~���W��q ~ q ~�t 2058ppw@$      sq ~���W��q ~ q ~�t 2059ppw@$      sq ~��~'�q ~ q ~�t 206ppw@$      sq ~���W�Iq ~ q ~�t 2060ppw@$      sq ~���W�
q ~ q ~�t 2061ppw@$      sq ~���W��q ~ q ~�t 2062ppw@$      sq ~���W��q ~ q ~�t 2063ppw@$      sq ~���W�Mq ~ q ~�t 2064ppw@$      sq ~���W�q ~ q ~�t 2065ppw@$      sq ~���X�q ~ q ~�t 2066ppw@$      sq ~���X�q ~ q ~�t 2067ppw@$      sq ~���X	Qq ~ q ~�t 2068ppw@$      sq ~���Xq ~ q ~�t 2069ppw@%_- ��sq ~��~+Jq ~ q ~�t 207ppw@$      sq ~���X_�q ~ q ~�t 2070ppw@$      sq ~���Xciq ~ q ~�t 2071ppw@$      sq ~���Xg*q ~ q ~�t 2072ppw@$      sq ~���Xj�q ~ q ~�t 2073ppw@$      sq ~���Xn�q ~ q ~�t 2074ppw@$      sq ~���Xrmq ~ q ~�t 2075ppw@$      sq ~���Xv.q ~ q ~�t 2076ppw@$      sq ~���Xy�q ~ q ~�t 2077ppw@$      sq ~���X}�q ~ q ~�t 2078ppw@$      sq ~���X�qq ~ q ~�t 2079ppw@$      sq ~��~/q ~ q ~�t 208ppw@$      sq ~���X�q ~ q ~�t 2080ppw@$      sq ~���X��q ~ q ~�t 2081ppw@$      sq ~���Xۉq ~ q ~�t 2082ppw@$      sq ~���X�Jq ~ q ~�t 2083ppw@$      sq ~���X�q ~ q ~�t 2084ppw@$      sq ~���X��q ~ q ~�t 2085ppw@$      sq ~���X�q ~ q ~�t 2086ppw@$      sq ~���X�Nq ~ q ~�t 2087ppw@$      sq ~���X�q ~ q ~�t 2088ppw@$      sq ~���X��q ~ q ~�t 2089ppw@$      sq ~��~2�q ~ q ~�t 209ppw@$      sq ~���YHfq ~ q ~�t 2090ppw@$      sq ~���YL'q ~ q ~�t 2091ppw@$      sq ~���YO�q ~ q ~�t 2092ppw@$      sq ~���YS�q ~ q ~�t 2093ppw@$      sq ~���YWjq ~ q ~�t 2094ppw@$      sq ~���Y[+q ~ q ~�t 2095ppw@$      sq ~���Y^�q ~ q ~�t 2096ppw@$      sq ~���Yb�q ~ q ~�t 2097ppw@%��_sq ~���Yfnq ~ q ~�t 2098ppw@$      sq ~���Yj/q ~ q ~�t 2099ppw@$      sq ~��{_fPq ~ q ~�t 21ppw@$      sq ~��~�bq ~ q ~�t 210ppw@$      sq ~���cH�q ~ q ~�t 2100ppw@$      sq ~���cLQq ~ q ~�t 2101ppw@$      sq ~���cPq ~ q ~�t 2102ppw@$      sq ~���cS�q ~ q ~�t 2103ppw@$      sq ~���cW�q ~ q ~�t 2104ppw@$      sq ~���c[Uq ~ q ~�t 2105ppw@$      sq ~���c_q ~ q ~�t 2106ppw@$      sq ~���cb�q ~ q ~�t 2107ppw@$      sq ~���cf�q ~ q ~�t 2108ppw@$      sq ~���cjYq ~ q ~�t 2109ppw@$      sq ~��~�#q ~ q ~�t 211ppw@$      sq ~���c��q ~ q ~�t 2110ppw@$      sq ~���c��q ~ q ~�t 2111ppw@$      sq ~���c�qq ~ q ~�t 2112ppw@$      sq ~���c�2q ~ q ~�t 2113ppw@$      sq ~���c��q ~ q ~�t 2114ppw@$      sq ~���cϴq ~ q ~�t 2115ppw@$      sq ~���c�uq ~ q ~�t 2116ppw@$      sq ~���c�6q ~ q ~�t 2117ppw@$      sq ~���c��q ~ q ~�t 2118ppw@$      sq ~���c޸q ~ q ~�t 2119ppw@$      sq ~��~��q ~ q ~�t 212ppw@
F[ sq ~���d1Nq ~ q ~�t 2120ppw@$      sq ~���d5q ~ q ~�t 2121ppw@$      sq ~���d8�q ~ q ~�t 2122ppw@$      sq ~���d<�q ~ q ~�t 2123ppw@$      sq ~���d@Rq ~ q ~�t 2124ppw@$      sq ~���dDq ~ q ~�t 2125ppw@$      sq ~���dG�q ~ q ~�t 2126ppw@%�e�_csq ~���dK�q ~ q ~�t 2127ppw@$      sq ~���dOVq ~ q ~�t 2128ppw@$      sq ~���dSq ~ q ~�t 2129ppw@$      sq ~��~��q ~ q ~�t 213ppw@$      sq ~���d��q ~ q ~�t 2130ppw@$      sq ~���d�nq ~ q ~�t 2131ppw@$      sq ~���d�/q ~ q ~�t 2132ppw@#�F��Fsq ~���d��q ~ q ~�t 2133ppw@$      sq ~���d��q ~ q ~�t 2134ppw@$      sq ~���d�rq ~ q ~�t 2135ppw@$      sq ~���d�3q ~ q ~�t 2136ppw@$      sq ~���d��q ~ q ~�t 2137ppw@$      sq ~���dõq ~ q ~�t 2138ppw@$      sq ~���d�vq ~ q ~�t 2139ppw@$      sq ~��~�fq ~ q ~�t 214ppw@$      sq ~���eq ~ q ~�t 2140ppw@$      sq ~���e�q ~ q ~�t 2141ppw@$      sq ~���e!�q ~ q ~�t 2142ppw@$      sq ~���e%Oq ~ q ~�t 2143ppw@ � ��'�sq ~���e)q ~ q ~�t 2144ppw@$      sq ~���e,�q ~ q ~�t 2145ppw@$      sq ~���e0�q ~ q ~�t 2146ppw@$      sq ~���e4Sq ~ q ~�t 2147ppw@$      sq ~���e8q ~ q ~�t 2148ppw@%�ʈ�Nsq ~���e;�q ~ q ~�t 2149ppw@$      sq ~��~�'q ~ q ~�t 215ppw@$      sq ~���e�kq ~ q ~�t 2150ppw@$      sq ~���e�,q ~ q ~�t 2151ppw@$      sq ~���e��q ~ q ~�t 2152ppw@$      sq ~���e��q ~ q ~�t 2153ppw@$      sq ~���e�oq ~ q ~�t 2154ppw@$      sq ~���e�0q ~ q ~�t 2155ppw@$      sq ~���e��q ~ q ~�t 2156ppw@$      sq ~���e��q ~ q ~�t 2157ppw@$      sq ~���e�sq ~ q ~�t 2158ppw@$      sq ~���e�4q ~ q ~�t 2159ppw@$      sq ~��~��q ~ q ~�t 216ppw@$      sq ~���f�q ~ q ~�t 2160ppw@$      sq ~���f�q ~ q ~�t 2161ppw@$      sq ~���f
Lq ~ q ~�t 2162ppw@$      sq ~���fq ~ q ~�t 2163ppw@$      sq ~���f�q ~ q ~�t 2164ppw@$      sq ~���f�q ~ q ~�t 2165ppw@$      sq ~���fPq ~ q ~�t 2166ppw@$      sq ~���fq ~ q ~�t 2167ppw@$      sq ~���f �q ~ q ~�t 2168ppw@$      sq ~���f$�q ~ q ~�t 2169ppw@$      sq ~��~��q ~ q ~�t 217ppw@$      sq ~���fw)q ~ q ~�t 2170ppw@$      sq ~���fz�q ~ q ~�t 2171ppw@$      sq ~���f~�q ~ q ~�t 2172ppw@$      sq ~���f�lq ~ q ~�t 2173ppw@$      sq ~���f�-q ~ q ~�t 2174ppw@$      sq ~���f��q ~ q ~�t 2175ppw@$      sq ~���f��q ~ q ~�t 2176ppw@$      sq ~���f�pq ~ q ~�t 2177ppw@$      sq ~���f�1q ~ q ~�t 2178ppw@$      sq ~���f��q ~ q ~�t 2179ppw@$      sq ~��~�jq ~ q ~�t 218ppw@$      sq ~���f�q ~ q ~�t 2180ppw@$      sq ~���f�Iq ~ q ~�t 2181ppw@$      sq ~���f�
q ~ q ~�t 2182ppw@$      sq ~���f��q ~ q ~�t 2183ppw@$      sq ~���f��q ~ q ~�t 2184ppw@$      sq ~���f�Mq ~ q ~�t 2185ppw@$      sq ~���gq ~ q ~�t 2186ppw@$      sq ~���g�q ~ q ~�t 2187ppw@$      sq ~���g	�q ~ q ~�t 2188ppw@$      sq ~���gQq ~ q ~�t 2189ppw@$      sq ~��~�+q ~ q ~�t 219ppw@$      sq ~���g_�q ~ q ~�t 2190ppw@$      sq ~���gc�q ~ q ~�t 2191ppw@$      sq ~���ggiq ~ q ~�t 2192ppw@$      sq ~���gk*q ~ q ~�t 2193ppw@$      sq ~���gn�q ~ q ~�t 2194ppw@$      sq ~���gr�q ~ q ~�t 2195ppw@$      sq ~���gvmq ~ q ~�t 2196ppw@$      sq ~���gz.q ~ q ~�t 2197ppw@$      sq ~���g}�q ~ q ~�t 2198ppw@*�E����sq ~���g��q ~ q ~�t 2199ppw@$      sq ~��{_jq ~ q ~�t 22ppw@3Mr�?csq ~��~��q ~ q ~�t 220ppw@$      sq ~���q`q ~ q ~�t 2200ppw@$      sq ~���qc�q ~ q ~�t 2201ppw@$      sq ~���qg�q ~ q ~�t 2202ppw@$      sq ~���qkTq ~ q ~�t 2203ppw@$      sq ~���qoq ~ q ~�t 2204ppw@$      sq ~���qr�q ~ q ~�t 2205ppw@$      sq ~���qv�q ~ q ~�t 2206ppw@$      sq ~���qzXq ~ q ~�t 2207ppw@$      sq ~���q~q ~ q ~�t 2208ppw@%ֆ"�ҵsq ~���q��q ~ q ~�t 2209ppw@$      sq ~��~��q ~ q ~�t 221ppw@$      sq ~���q�pq ~ q ~�t 2210ppw@$      sq ~���q�1q ~ q ~�t 2211ppw@$      sq ~���q��q ~ q ~�t 2212ppw@#�hr�Nsq ~���q߳q ~ q ~�t 2213ppw@$      sq ~���q�tq ~ q ~�t 2214ppw@$      sq ~���q�5q ~ q ~�t 2215ppw@$      sq ~���q��q ~ q ~�t 2216ppw@$      sq ~���q�q ~ q ~�t 2217ppw@$      sq ~���q�xq ~ q ~�t 2218ppw@$      sq ~���q�9q ~ q ~�t 2219ppw@$      sq ~��~ Cq ~ q ~�t 222ppw@$      sq ~���rH�q ~ q ~�t 2220ppw@$      sq ~���rL�q ~ q ~�t 2221ppw@$      sq ~���rPQq ~ q ~�t 2222ppw@$      sq ~���rTq ~ q ~�t 2223ppw@$      sq ~���rW�q ~ q ~�t 2224ppw@$      sq ~���r[�q ~ q ~�t 2225ppw@$      sq ~���r_Uq ~ q ~�t 2226ppw@$      sq ~���rcq ~ q ~�t 2227ppw@$      sq ~���rf�q ~ q ~�t 2228ppw@$      sq ~���rj�q ~ q ~�t 2229ppw@$      sq ~��~ q ~ q ~�t 223ppw@$      sq ~���r�.q ~ q ~�t 2230ppw@$      sq ~���r��q ~ q ~�t 2231ppw@$      sq ~���rİq ~ q ~�t 2232ppw@$      sq ~���r�qq ~ q ~�t 2233ppw@$      sq ~���r�2q ~ q ~�t 2234ppw@$      sq ~���r��q ~ q ~�t 2235ppw@$      sq ~���rӴq ~ q ~�t 2236ppw@$      sq ~���r�uq ~ q ~�t 2237ppw@$      sq ~���r�6q ~ q ~�t 2238ppw@$      sq ~���r��q ~ q ~�t 2239ppw@$      sq ~��~ �q ~ q ~�t 224ppw@$      sq ~���s1�q ~ q ~�t 2240ppw@$      sq ~���s5Nq ~ q ~�t 2241ppw@$      sq ~���s9q ~ q ~�t 2242ppw@$      sq ~���s<�q ~ q ~�t 2243ppw@$      sq ~���s@�q ~ q ~�t 2244ppw@$      sq ~���sDRq ~ q ~�t 2245ppw@$      sq ~���sHq ~ q ~�t 2246ppw@$      sq ~���sK�q ~ q ~�t 2247ppw@$      sq ~���sO�q ~ q ~�t 2248ppw@$      sq ~���sSVq ~ q ~�t 2249ppw@$      sq ~��~ �q ~ q ~�t 225ppw@$      sq ~���s��q ~ q ~�t 2250ppw@$      sq ~���s��q ~ q ~�t 2251ppw@$      sq ~���s�nq ~ q ~�t 2252ppw@$      sq ~���s�/q ~ q ~�t 2253ppw@$      sq ~���s��q ~ q ~�t 2254ppw@$      sq ~���s��q ~ q ~�t 2255ppw@$      sq ~���s�rq ~ q ~�t 2256ppw@$      sq ~���s�3q ~ q ~�t 2257ppw@$      sq ~���s��q ~ q ~�t 2258ppw@$      sq ~���sǵq ~ q ~�t 2259ppw@$      sq ~��~ Gq ~ q ~�t 226ppw@$      sq ~���tKq ~ q ~�t 2260ppw@$      sq ~���tq ~ q ~�t 2261ppw@$      sq ~���t!�q ~ q ~�t 2262ppw@'�����sq ~���t%�q ~ q ~�t 2263ppw@$      sq ~���t)Oq ~ q ~�t 2264ppw@$      sq ~���t-q ~ q ~�t 2265ppw@$      sq ~���t0�q ~ q ~�t 2266ppw@%��� ��sq ~���t4�q ~ q ~�t 2267ppw@$      sq ~���t8Sq ~ q ~�t 2268ppw@$      sq ~���t<q ~ q ~�t 2269ppw@$      sq ~��~ q ~ q ~�t 227ppw@$      sq ~���t��q ~ q ~�t 2270ppw@$      sq ~���t�kq ~ q ~�t 2271ppw@$      sq ~���t�,q ~ q ~�t 2272ppw@$      sq ~���t��q ~ q ~�t 2273ppw@$      sq ~���t��q ~ q ~�t 2274ppw@$      sq ~���t�oq ~ q ~�t 2275ppw@$      sq ~���t�0q ~ q ~�t 2276ppw@$      sq ~���t��q ~ q ~�t 2277ppw@$      sq ~���t��q ~ q ~�t 2278ppw@$      sq ~���t�sq ~ q ~�t 2279ppw@$      sq ~��~ �q ~ q ~�t 228ppw@$      sq ~���u	q ~ q ~�t 2280ppw@$      sq ~���u�q ~ q ~�t 2281ppw@$      sq ~���u
�q ~ q ~�t 2282ppw@$      sq ~���uLq ~ q ~�t 2283ppw@$      sq ~���uq ~ q ~�t 2284ppw@$      sq ~���u�q ~ q ~�t 2285ppw@$      sq ~���u�q ~ q ~�t 2286ppw@$      sq ~���uPq ~ q ~�t 2287ppw@$      sq ~���u!q ~ q ~�t 2288ppw@$      sq ~���u$�q ~ q ~�t 2289ppw@$      sq ~��~ �q ~ q ~�t 229ppw@$      sq ~���uwhq ~ q ~�t 2290ppw@$      sq ~���u{)q ~ q ~�t 2291ppw@$      sq ~���u~�q ~ q ~�t 2292ppw@$      sq ~���u��q ~ q ~�t 2293ppw@$      sq ~���u�lq ~ q ~�t 2294ppw@$      sq ~���u�-q ~ q ~�t 2295ppw@$      sq ~���u��q ~ q ~�t 2296ppw@$      sq ~���u��q ~ q ~�t 2297ppw@$      sq ~���u�pq ~ q ~�t 2298ppw@$      sq ~���u�1q ~ q ~�t 2299ppw@$      sq ~��{_m�q ~ q ~�t 23ppw@%�]���ssq ~��~ n q ~ q ~�t 230ppw@$      sq ~���w�q ~ q ~�t 2300ppw@$      sq ~���{Sq ~ q ~�t 2301ppw@$      sq ~���q ~ q ~�t 2302ppw@$      sq ~�����q ~ q ~�t 2303ppw@$      sq ~�����q ~ q ~�t 2304ppw@$      sq ~����Wq ~ q ~�t 2305ppw@$      sq ~����q ~ q ~�t 2306ppw@$      sq ~�����q ~ q ~�t 2307ppw@$      sq ~�����q ~ q ~�t 2308ppw@$      sq ~����[q ~ q ~�t 2309ppw@$      sq ~��~ q�q ~ q ~�t 231ppw@$      sq ~�����q ~ q ~�t 2310ppw@$      sq ~����q ~ q ~�t 2311ppw@$      sq ~����sq ~ q ~�t 2312ppw@$      sq ~����4q ~ q ~�t 2313ppw@$      sq ~�����q ~ q ~�t 2314ppw@$      sq ~�����q ~ q ~�t 2315ppw@$      sq ~��Ӏwq ~ q ~�t 2316ppw@$      sq ~��Ӏ8q ~ q ~�t 2317ppw@$      sq ~��Ӏ	�q ~ q ~�t 2318ppw@$      sq ~��Ӏ�q ~ q ~�t 2319ppw@$      sq ~��~ u�q ~ q ~�t 232ppw@$      sq ~��Ӏ`Pq ~ q ~�t 2320ppw@$      sq ~��Ӏdq ~ q ~�t 2321ppw@$      sq ~��Ӏg�q ~ q ~�t 2322ppw@$      sq ~��Ӏk�q ~ q ~�t 2323ppw@$      sq ~��ӀoTq ~ q ~�t 2324ppw@$      sq ~��Ӏsq ~ q ~�t 2325ppw@$      sq ~��Ӏv�q ~ q ~�t 2326ppw@$      sq ~��Ӏz�q ~ q ~�t 2327ppw@$      sq ~��Ӏ~Xq ~ q ~�t 2328ppw@$7��O�sq ~��Ӏ�q ~ q ~�t 2329ppw@$      sq ~��~ ycq ~ q ~�t 233ppw@$      sq ~��Ӏԯq ~ q ~�t 2330ppw@$      sq ~��Ӏ�pq ~ q ~�t 2331ppw@$      sq ~��Ӏ�1q ~ q ~�t 2332ppw@$      sq ~��Ӏ��q ~ q ~�t 2333ppw@$      sq ~��Ӏ�q ~ q ~�t 2334ppw@$      sq ~��Ӏ�tq ~ q ~�t 2335ppw@$      sq ~��Ӏ�5q ~ q ~�t 2336ppw@$      sq ~��Ӏ��q ~ q ~�t 2337ppw@$      sq ~��Ӏ�q ~ q ~�t 2338ppw@$      sq ~��Ӏ�xq ~ q ~�t 2339ppw@$      sq ~��~ }$q ~ q ~�t 234ppw@$      sq ~��ӁIq ~ q ~�t 2340ppw@$      sq ~��ӁL�q ~ q ~�t 2341ppw@$      sq ~��ӁP�q ~ q ~�t 2342ppw@$      sq ~��ӁTQq ~ q ~�t 2343ppw@$      sq ~��ӁXq ~ q ~�t 2344ppw@$      sq ~��Ӂ[�q ~ q ~�t 2345ppw@$      sq ~��Ӂ_�q ~ q ~�t 2346ppw@$      sq ~��ӁcUq ~ q ~�t 2347ppw@$      sq ~��Ӂgq ~ q ~�t 2348ppw@$      sq ~��Ӂj�q ~ q ~�t 2349ppw@$      sq ~��~ ��q ~ q ~�t 235ppw@$      sq ~��Ӂ�mq ~ q ~�t 2350ppw@$      sq ~��Ӂ�.q ~ q ~�t 2351ppw@$      sq ~��Ӂ��q ~ q ~�t 2352ppw@$      sq ~��ӁȰq ~ q ~�t 2353ppw@$      sq ~��Ӂ�qq ~ q ~�t 2354ppw@$      sq ~��Ӂ�2q ~ q ~�t 2355ppw@$      sq ~��Ӂ��q ~ q ~�t 2356ppw@$      sq ~��Ӂ״q ~ q ~�t 2357ppw@$      sq ~��Ӂ�uq ~ q ~�t 2358ppw@$      sq ~��Ӂ�6q ~ q ~�t 2359ppw@$      sq ~��~ ��q ~ q ~�t 236ppw@$      sq ~��ӂ1�q ~ q ~�t 2360ppw@$      sq ~��ӂ5�q ~ q ~�t 2361ppw@$      sq ~��ӂ9Nq ~ q ~�t 2362ppw@$      sq ~��ӂ=q ~ q ~�t 2363ppw@$      sq ~��ӂ@�q ~ q ~�t 2364ppw@$      sq ~��ӂD�q ~ q ~�t 2365ppw@$      sq ~��ӂHRq ~ q ~�t 2366ppw@$      sq ~��ӂLq ~ q ~�t 2367ppw@$      sq ~��ӂO�q ~ q ~�t 2368ppw@$      sq ~��ӂS�q ~ q ~�t 2369ppw@$      sq ~��~ �gq ~ q ~�t 237ppw@$      sq ~��ӂ�+q ~ q ~�t 2370ppw@$      sq ~��ӂ��q ~ q ~�t 2371ppw@$      sq ~��ӂ��q ~ q ~�t 2372ppw@$      sq ~��ӂ�nq ~ q ~�t 2373ppw@$      sq ~��ӂ�/q ~ q ~�t 2374ppw@$      sq ~��ӂ��q ~ q ~�t 2375ppw@$      sq ~��ӂ��q ~ q ~�t 2376ppw@$      sq ~��ӂ�rq ~ q ~�t 2377ppw@$      sq ~��ӂ�3q ~ q ~�t 2378ppw@$      sq ~��ӂ��q ~ q ~�t 2379ppw@$      sq ~��~ �(q ~ q ~�t 238ppw@$      sq ~��Ӄ�q ~ q ~�t 2380ppw@$      sq ~��ӃKq ~ q ~�t 2381ppw@#��o�"sq ~��Ӄ"q ~ q ~�t 2382ppw@$      sq ~��Ӄ%�q ~ q ~�t 2383ppw@$      sq ~��Ӄ)�q ~ q ~�t 2384ppw@$      sq ~��Ӄ-Oq ~ q ~�t 2385ppw@$      sq ~��Ӄ1q ~ q ~�t 2386ppw@$      sq ~��Ӄ4�q ~ q ~�t 2387ppw@$      sq ~��Ӄ8�q ~ q ~�t 2388ppw@$      sq ~��Ӄ<Sq ~ q ~�t 2389ppw@$      sq ~��~ ��q ~ q ~�t 239ppw@$      sq ~��Ӄ��q ~ q ~�t 2390ppw@$      sq ~��Ӄ��q ~ q ~�t 2391ppw@$      sq ~��Ӄ�kq ~ q ~�t 2392ppw@$      sq ~��Ӄ�,q ~ q ~�t 2393ppw@$      sq ~��Ӄ��q ~ q ~�t 2394ppw@$      sq ~��Ӄ��q ~ q ~�t 2395ppw@$      sq ~��Ӄ�oq ~ q ~�t 2396ppw@%�/�ͭ>sq ~��Ӄ�0q ~ q ~�t 2397ppw@$      sq ~��Ӄ��q ~ q ~�t 2398ppw@$      sq ~��Ӄ��q ~ q ~�t 2399ppw@$      sq ~��{_q�q ~ q ~�t 24ppw@7�76�Rsq ~��~ �q ~ q ~�t 240ppw@$      sq ~��Ӎ�q ~ q ~�t 2400ppw@$      sq ~��Ӎ��q ~ q ~�t 2401ppw@$      sq ~��Ӎ��q ~ q ~�t 2402ppw@$      sq ~��Ӎ�Vq ~ q ~�t 2403ppw@$      sq ~��Ӎ�q ~ q ~�t 2404ppw@$      sq ~��Ӎ��q ~ q ~�t 2405ppw@$      sq ~��Ӎ��q ~ q ~�t 2406ppw@)�J
�sq ~��Ӎ�Zq ~ q ~�t 2407ppw@$      sq ~��Ӎ�q ~ q ~�t 2408ppw@$      sq ~��Ӎ��q ~ q ~�t 2409ppw@$      sq ~��~ �@q ~ q ~�t 241ppw@$      sq ~��ӎrq ~ q ~�t 2410ppw@$      sq ~��ӎ3q ~ q ~�t 2411ppw@$      sq ~��ӎ
�q ~ q ~�t 2412ppw@$      sq ~��ӎ�q ~ q ~�t 2413ppw@'L�L��sq ~��ӎvq ~ q ~�t 2414ppw@$      sq ~��ӎ7q ~ q ~�t 2415ppw@$      sq ~��ӎ�q ~ q ~�t 2416ppw@$      sq ~��ӎ�q ~ q ~�t 2417ppw@$      sq ~��ӎ!zq ~ q ~�t 2418ppw@$      sq ~��ӎ%;q ~ q ~�t 2419ppw@$      sq ~��~ �q ~ q ~�t 242ppw@$      sq ~��ӎw�q ~ q ~�t 2420ppw@$      sq ~��ӎ{�q ~ q ~�t 2421ppw@$      sq ~��ӎSq ~ q ~�t 2422ppw@$      sq ~��ӎ�q ~ q ~�t 2423ppw@$      sq ~��ӎ��q ~ q ~�t 2424ppw@$      sq ~��ӎ��q ~ q ~�t 2425ppw@$      sq ~��ӎ�Wq ~ q ~�t 2426ppw@$      sq ~��ӎ�q ~ q ~�t 2427ppw@$      sq ~��ӎ��q ~ q ~�t 2428ppw@$      sq ~��ӎ��q ~ q ~�t 2429ppw@%��Kߢ�sq ~��~ ��q ~ q ~�t 243ppw@$      sq ~��ӎ�0q ~ q ~�t 2430ppw@$      sq ~��ӎ��q ~ q ~�t 2431ppw@$      sq ~��ӎ�q ~ q ~�t 2432ppw@$      sq ~��ӎ�sq ~ q ~�t 2433ppw@$      sq ~��ӎ�4q ~ q ~�t 2434ppw@$      sq ~��ӎ��q ~ q ~�t 2435ppw@$      sq ~��ӏ�q ~ q ~�t 2436ppw@$      sq ~��ӏwq ~ q ~�t 2437ppw@$      sq ~��ӏ
8q ~ q ~�t 2438ppw@$      sq ~��ӏ�q ~ q ~�t 2439ppw@$      sq ~��~ �q ~ q ~�t 244ppw@$      sq ~��ӏ`�q ~ q ~�t 2440ppw@$      sq ~��ӏdPq ~ q ~�t 2441ppw@$      sq ~��ӏhq ~ q ~�t 2442ppw@$      sq ~��ӏk�q ~ q ~�t 2443ppw@$      sq ~��ӏo�q ~ q ~�t 2444ppw@$      sq ~��ӏsTq ~ q ~�t 2445ppw@$      sq ~��ӏwq ~ q ~�t 2446ppw@$      sq ~��ӏz�q ~ q ~�t 2447ppw@$      sq ~��ӏ~�q ~ q ~�t 2448ppw@$      sq ~��ӏ�Xq ~ q ~�t 2449ppw@$      sq ~��~ �Dq ~ q ~�t 245ppw@$      sq ~��ӏ��q ~ q ~�t 2450ppw@$      sq ~��ӏدq ~ q ~�t 2451ppw@$      sq ~��ӏ�pq ~ q ~�t 2452ppw@$      sq ~��ӏ�1q ~ q ~�t 2453ppw@$      sq ~��ӏ��q ~ q ~�t 2454ppw@$      sq ~��ӏ�q ~ q ~�t 2455ppw@$      sq ~��ӏ�tq ~ q ~�t 2456ppw@$      sq ~��ӏ�5q ~ q ~�t 2457ppw@$      sq ~��ӏ��q ~ q ~�t 2458ppw@$      sq ~��ӏ��q ~ q ~�t 2459ppw@&��]8�sq ~��~ �q ~ q ~�t 246ppw@$      sq ~��ӐIMq ~ q ~�t 2460ppw@$      sq ~��ӐMq ~ q ~�t 2461ppw@$      sq ~��ӐP�q ~ q ~�t 2462ppw@$      sq ~��ӐT�q ~ q ~�t 2463ppw@$      sq ~��ӐXQq ~ q ~�t 2464ppw@$      sq ~��Ӑ\q ~ q ~�t 2465ppw@$      sq ~��Ӑ_�q ~ q ~�t 2466ppw@$      sq ~��Ӑc�q ~ q ~�t 2467ppw@$      sq ~��ӐgUq ~ q ~�t 2468ppw@$      sq ~��Ӑkq ~ q ~�t 2469ppw@$      sq ~��~ ��q ~ q ~�t 247ppw@$      sq ~��Ӑ��q ~ q ~�t 2470ppw@$      sq ~��Ӑ�mq ~ q ~�t 2471ppw@%����\sq ~��Ӑ�.q ~ q ~�t 2472ppw@$      sq ~��Ӑ��q ~ q ~�t 2473ppw@$      sq ~��Ӑ̰q ~ q ~�t 2474ppw@$      sq ~��Ӑ�qq ~ q ~�t 2475ppw@$      sq ~��Ӑ�2q ~ q ~�t 2476ppw@$      sq ~��Ӑ��q ~ q ~�t 2477ppw@$      sq ~��Ӑ۴q ~ q ~�t 2478ppw@$      sq ~��Ӑ�uq ~ q ~�t 2479ppw@$      sq ~��~! �q ~ q ~�t 248ppw@$      sq ~��ӑ2q ~ q ~�t 2480ppw@$      sq ~��ӑ5�q ~ q ~�t 2481ppw@$      sq ~��ӑ9�q ~ q ~�t 2482ppw@$      sq ~��ӑ=Nq ~ q ~�t 2483ppw@$      sq ~��ӑAq ~ q ~�t 2484ppw@$      sq ~��ӑD�q ~ q ~�t 2485ppw@$      sq ~��ӑH�q ~ q ~�t 2486ppw?�      sq ~��ӑLRq ~ q ~�t 2487ppw?��.NF�(sq ~��ӑPq ~ q ~�t 2488ppw@O��k#5sq ~��ӑS�q ~ q ~�t 2489ppw?������sq ~��~!Hq ~ q ~�t 249ppw@$      sq ~��ӑ�jq ~ q ~�t 2490ppw@��躟�sq ~��ӑ�+q ~ q ~�t 2491ppw@�X�S3sq ~��ӑ��q ~ q ~�t 2492ppw?��E>�Ysq ~��ӑ��q ~ q ~�t 2493ppw@ �
F��sq ~��ӑ�nq ~ q ~�t 2494ppw?��s���sq ~��ӑ�/q ~ q ~�t 2495ppw@!�$�!|sq ~��ӑ��q ~ q ~�t 2496ppw@���?�sq ~��ӑ��q ~ q ~�t 2497ppw��̂�tsq ~��ӑ�rq ~ q ~�t 2498ppw�Н�ޝ�sq ~��ӑ�3q ~ q ~�t 2499ppw@,�
�g��sq ~��{_uTq ~ q ~�t 25ppw@$      sq ~��~!V�q ~ q ~�t 250ppw@$      sq ~��ӛ��q ~ q ~�t 2500ppw?�SH�SVsq ~��ӛ�Uq ~ q ~�t 2501ppw?�L��Ҿ/sq ~��ӛ�q ~ q ~�t 2502ppw@�����5sq ~��ӛ��q ~ q ~�t 2503ppw?��G��sq ~��ӛ��q ~ q ~�t 2504ppw?�@�`e��sq ~��ӛ�Yq ~ q ~�t 2505ppw?�@�`e��sq ~��ӛ�q ~ q ~�t 2506ppw?�@�`e��sq ~��ӛ��q ~ q ~�t 2507ppw?�@�`e��sq ~��ӛĜq ~ q ~�t 2508ppw?�@�`e��sq ~��ӛ�]q ~ q ~�t 2509ppw?�Xs��^sq ~��~!Z�q ~ q ~�t 251ppw@$      sq ~��Ӝ�q ~ q ~�t 2510ppw?����#�sq ~��Ӝ�q ~ q ~�t 2511ppw@#���!Rsq ~��Ӝ"uq ~ q ~�t 2512ppw?���5�V�sq ~��Ӝ&6q ~ q ~�t 2513ppw?��b�ȟ�sq ~��Ӝ)�q ~ q ~�t 2514ppw@�����7sq ~��Ӝ-�q ~ q ~�t 2515ppw?�� ^��sq ~��Ӝ1yq ~ q ~�t 2516ppw?�����h_sq ~��Ӝ5:q ~ q ~�t 2517ppw@�!�j�sq ~��Ӝ8�q ~ q ~�t 2518ppw?��O�b8�sq ~��Ӝ<�q ~ q ~�t 2519ppw@�GD��sq ~��~!^`q ~ q ~�t 252ppw@$      sq ~��Ӝ�Rq ~ q ~�t 2520ppw?�/73�sq ~��Ӝ�q ~ q ~�t 2521ppw?��\�h�sq ~��Ӝ��q ~ q ~�t 2522ppw�,pP*]�sq ~��Ӝ��q ~ q ~�t 2523ppw?����sq ~��Ӝ�Vq ~ q ~�t 2524ppw?��=��sq ~��Ӝ�q ~ q ~�t 2525ppw?��=��sq ~��Ӝ��q ~ q ~�t 2526ppw?���$Kfsq ~��Ӝ��q ~ q ~�t 2527ppw?�����G3sq ~��Ӝ�Zq ~ q ~�t 2528ppw?�����O+sq ~��Ӝ�q ~ q ~�t 2529ppw?�ݼ���Nsq ~��~!b!q ~ q ~�t 253ppw@$      sq ~��ӝ�q ~ q ~�t 2530ppw?��M�*Osq ~��ӝrq ~ q ~�t 2531ppw?��M�*Osq ~��ӝ3q ~ q ~�t 2532ppw?��x��bsq ~��ӝ�q ~ q ~�t 2533ppw?�EӪ�n{sq ~��ӝ�q ~ q ~�t 2534ppw����\��sq ~��ӝvq ~ q ~�t 2535ppw@"�͞�y*sq ~��ӝ7q ~ q ~�t 2536ppw@Ʋ'�)�sq ~��ӝ�q ~ q ~�t 2537ppw?��0�~��sq ~��ӝ!�q ~ q ~�t 2538ppw?�[C_�j�sq ~��ӝ%zq ~ q ~�t 2539ppw?�[C_�j�sq ~��~!e�q ~ q ~�t 254ppw@$      sq ~��ӝxq ~ q ~�t 2540ppw?��0�~��sq ~��ӝ{�q ~ q ~�t 2541ppw@��=��Zsq ~��ӝ�q ~ q ~�t 2542ppw@%�{^m��sq ~��ӝ�Sq ~ q ~�t 2543ppw@�<픃xsq ~��ӝ�q ~ q ~�t 2544ppw@$#�Ю�sq ~��ӝ��q ~ q ~�t 2545ppw?�e
�`��sq ~��ӝ��q ~ q ~�t 2546ppw?�����sq ~��ӝ�Wq ~ q ~�t 2547ppw?�<�Ǯ�ksq ~��ӝ�q ~ q ~�t 2548ppw?０���sq ~��ӝ��q ~ q ~�t 2549ppw?�X$W��sq ~��~!i�q ~ q ~�t 255ppw@$      sq ~��ӝ�oq ~ q ~�t 2550ppw@^��&Msq ~��ӝ�0q ~ q ~�t 2551ppw���xRhsq ~��ӝ��q ~ q ~�t 2552ppw@�Q��sq ~��ӝ��q ~ q ~�t 2553ppw@�/شsq ~��ӝ�sq ~ q ~�t 2554ppw?�A�&�sq ~��ӝ�4q ~ q ~�t 2555ppw?�qWk�wsq ~��Ӟ�q ~ q ~�t 2556ppw?�A�$�sq ~��Ӟ�q ~ q ~�t 2557ppw� �K ��sq ~��Ӟ
wq ~ q ~�t 2558ppw?ΡO�ybRsq ~��Ӟ8q ~ q ~�t 2559ppw?�%ԩ��sq ~��~!mdq ~ q ~�t 256ppw@$      sq ~��Ӟ`�q ~ q ~�t 2560ppw?��2O�*psq ~��Ӟd�q ~ q ~�t 2561ppw?�%ԩ��sq ~��ӞhPq ~ q ~�t 2562ppw?�cy�q9\sq ~��Ӟlq ~ q ~�t 2563ppw?�eDa��sq ~��Ӟo�q ~ q ~�t 2564ppw?�q;.6$sq ~��Ӟs�q ~ q ~�t 2565ppw?��U��6�sq ~��ӞwTq ~ q ~�t 2566ppw���f#,��sq ~��Ӟ{q ~ q ~�t 2567ppw?9�sq ~��Ӟ~�q ~ q ~�t 2568ppw?��=��sq ~��Ӟ��q ~ q ~�t 2569ppw?���v�sq ~��~!q%q ~ q ~�t 257ppw@$      sq ~��Ӟ�-q ~ q ~�t 2570ppw?���v�sq ~��Ӟ��q ~ q ~�t 2571ppw?��+�;
sq ~��Ӟܯq ~ q ~�t 2572ppw@
` ��sq ~��Ӟ�pq ~ q ~�t 2573ppw?�|�����sq ~��Ӟ�1q ~ q ~�t 2574ppw���I���sq ~��Ӟ��q ~ q ~�t 2575ppw@#�r�͚sq ~��Ӟ�q ~ q ~�t 2576ppw@_S��7Dsq ~��Ӟ�tq ~ q ~�t 2577ppw?�o&�$�sq ~��Ӟ�5q ~ q ~�t 2578ppw?�m���sq ~��Ӟ��q ~ q ~�t 2579ppw?�jiAKV�sq ~��~!t�q ~ q ~�t 258ppw@$      sq ~��ӟI�q ~ q ~�t 2580ppw?�h]sq ~��ӟMMq ~ q ~�t 2581ppw?�h]sq ~��ӟQq ~ q ~�t 2582ppw@6���sq ~��ӟT�q ~ q ~�t 2583ppw@oY,�sq ~��ӟX�q ~ q ~�t 2584ppw?�=��"�`sq ~��ӟ\Qq ~ q ~�t 2585ppw?�=��"��sq ~��ӟ`q ~ q ~�t 2586ppw��)�6=�sq ~��ӟc�q ~ q ~�t 2587ppw?�Y�Gsq ~��ӟg�q ~ q ~�t 2588ppw?�XJӗ2�sq ~��ӟkUq ~ q ~�t 2589ppw?�S�<��sq ~��~!x�q ~ q ~�t 259ppw@$      sq ~��ӟ��q ~ q ~�t 2590ppw?���H?sq ~��ӟ��q ~ q ~�t 2591ppw���8���sq ~��ӟ�mq ~ q ~�t 2592ppw?���o�-Esq ~��ӟ�.q ~ q ~�t 2593ppw?�K�f�}vsq ~��ӟ��q ~ q ~�t 2594ppw@Ô�	Rsq ~��ӟаq ~ q ~�t 2595ppw��E&���sq ~��ӟ�qq ~ q ~�t 2596ppw@��8�
sq ~��ӟ�2q ~ q ~�t 2597ppw?�G�1$sq ~��ӟ��q ~ q ~�t 2598ppw?�BX-b4sq ~��ӟߴq ~ q ~�t 2599ppw?�<�O��sq ~��{_yq ~ q ~�t 26ppw@T16���sq ~��~!�=q ~ q ~�t 260ppw@$      sq ~��ө�q ~ q ~�t 2600ppw?�5�K�#sq ~��ө��q ~ q ~�t 2601ppw?�4LcZ��sq ~��өŗq ~ q ~�t 2602ppw?�4LcZ�usq ~��ө�Xq ~ q ~�t 2603ppw?�4LcZ�usq ~��ө�q ~ q ~�t 2604ppw?�{�B���sq ~��ө��q ~ q ~�t 2605ppw?�.O��sq ~��өԛq ~ q ~�t 2606ppw@֨K��sq ~��ө�\q ~ q ~�t 2607ppw?�c�����sq ~��ө�q ~ q ~�t 2608ppw        sq ~��ө��q ~ q ~�t 2609ppw        sq ~��~!��q ~ q ~�t 261ppw@$      sq ~��Ӫ2tq ~ q ~�t 2610ppw?���W-"sq ~��Ӫ65q ~ q ~�t 2611ppw?�Z���|sq ~��Ӫ9�q ~ q ~�t 2612ppw?��>�e sq ~��Ӫ=�q ~ q ~�t 2613ppw?�5�x���sq ~��ӪAxq ~ q ~�t 2614ppw?�J�I_sq ~��ӪE9q ~ q ~�t 2615ppw?����sq ~��ӪH�q ~ q ~�t 2616ppw?��lp��sq ~��ӪL�q ~ q ~�t 2617ppw?��U��sq ~��ӪP|q ~ q ~�t 2618ppw?���O Zsq ~��ӪT=q ~ q ~�t 2619ppw?��b8sq ~��~!ҿq ~ q ~�t 262ppw@$      sq ~��Ӫ��q ~ q ~�t 2620ppw?�ϊyÏ�sq ~��Ӫ��q ~ q ~�t 2621ppw?���+RJsq ~��Ӫ�Uq ~ q ~�t 2622ppw?޿��W[�sq ~��Ӫ�q ~ q ~�t 2623ppw?޿��W[�sq ~��Ӫ��q ~ q ~�t 2624ppw?�Չ�K�sq ~��Ӫ��q ~ q ~�t 2625ppw?�[<?�Xsq ~��Ӫ�Yq ~ q ~�t 2626ppw?��DsE}sq ~��Ӫ�q ~ q ~�t 2627ppw@@˜�	sq ~��Ӫ��q ~ q ~�t 2628ppw?�K�sq ~��ӪȜq ~ q ~�t 2629ppw?��G11��sq ~��~!րq ~ q ~�t 263ppw@$      sq ~��ӫ2q ~ q ~�t 2630ppw@�c{Ĕsq ~��ӫ�q ~ q ~�t 2631ppw��0-w�1@sq ~��ӫ"�q ~ q ~�t 2632ppw@��m��
sq ~��ӫ&uq ~ q ~�t 2633ppw@���sq ~��ӫ*6q ~ q ~�t 2634ppw?���.�sq ~��ӫ-�q ~ q ~�t 2635ppw?�<՛sq ~��ӫ1�q ~ q ~�t 2636ppw?��$l��sq ~��ӫ5yq ~ q ~�t 2637ppw?��4p!sq ~��ӫ9:q ~ q ~�t 2638ppw?����Ksq ~��ӫ<�q ~ q ~�t 2639ppw?���sq ~��~!�Aq ~ q ~�t 264ppw@$      sq ~��ӫ��q ~ q ~�t 2640ppw?�z���~�sq ~��ӫ�Rq ~ q ~�t 2641ppw?�v�	���sq ~��ӫ�q ~ q ~�t 2642ppw?�s��-vsq ~��ӫ��q ~ q ~�t 2643ppw?�s��-vsq ~��ӫ��q ~ q ~�t 2644ppw?�c�WG=wsq ~��ӫ�Vq ~ q ~�t 2645ppw@(��eJ�sq ~��ӫ�q ~ q ~�t 2646ppw�b�T��sq ~��ӫ��q ~ q ~�t 2647ppw?՚�d©sq ~��ӫ��q ~ q ~�t 2648ppw?�����sq ~��ӫ�Zq ~ q ~�t 2649ppw��D9��sq ~��~!�q ~ q ~�t 265ppw@$      sq ~��Ӭ�q ~ q ~�t 2650ppw?�N�����sq ~��Ӭ�q ~ q ~�t 2651ppw?�dߌ
1-sq ~��Ӭrq ~ q ~�t 2652ppw@
��z��sq ~��Ӭ3q ~ q ~�t 2653ppw@9�ɉ0sq ~��Ӭ�q ~ q ~�t 2654ppw?��e�+sq ~��Ӭ�q ~ q ~�t 2655ppw��Z{=�csq ~��Ӭvq ~ q ~�t 2656ppw        sq ~��~!��q ~ q ~�t 266ppw@$      sq ~��~!�q ~ q ~�t 267ppw@$      sq ~��~!�Eq ~ q ~�t 268ppw@$      sq ~��~!�q ~ q ~�t 269ppw@$      sq ~��{_|�q ~ q ~�t 27ppw@$      sq ~��~"?�q ~ q ~�t 270ppw@$      sq ~��~"C]q ~ q ~�t 271ppw@$      sq ~��~"Gq ~ q ~�t 272ppw@$      sq ~��~"J�q ~ q ~�t 273ppw@$      sq ~��~"N�q ~ q ~�t 274ppw@$      sq ~��~"Raq ~ q ~�t 275ppw@$      sq ~��~"V"q ~ q ~�t 276ppw@$      sq ~��~"Y�q ~ q ~�t 277ppw@$      sq ~��~"]�q ~ q ~�t 278ppw@$      sq ~��~"aeq ~ q ~�t 279ppw@$      sq ~��{_��q ~ q ~�t 28ppw@$      sq ~��~"��q ~ q ~�t 280ppw@$      sq ~��~"��q ~ q ~�t 281ppw@$      sq ~��~"�}q ~ q ~�t 282ppw@$      sq ~��~"�>q ~ q ~�t 283ppw@$      sq ~��~"��q ~ q ~�t 284ppw@$      sq ~��~"��q ~ q ~�t 285ppw@$      sq ~��~"ʁq ~ q ~�t 286ppw@$      sq ~��~"�Bq ~ q ~�t 287ppw@$      sq ~��~"�q ~ q ~�t 288ppw@$      sq ~��~"��q ~ q ~�t 289ppw@$      sq ~��{_�Xq ~ q ~�t 29ppw@+�Ք��sq ~��~#(Zq ~ q ~�t 290ppw@$      sq ~��~#,q ~ q ~�t 291ppw@$      sq ~��~#/�q ~ q ~�t 292ppw@$      sq ~��~#3�q ~ q ~�t 293ppw@$      sq ~��~#7^q ~ q ~�t 294ppw@$      sq ~��~#;q ~ q ~�t 295ppw@$      sq ~��~#>�q ~ q ~�t 296ppw@$      sq ~��~#B�q ~ q ~�t 297ppw@$      sq ~��~#Fbq ~ q ~�t 298ppw@$      sq ~��~#J#q ~ q ~�t 299ppw@$      sq ~��{H�Dq ~ q ~�t 3ppw@$      sq ~��{_��q ~ q ~�t 30ppw@$      sq ~��~-(�q ~ q ~�t 300ppw@$      sq ~��~-,Eq ~ q ~�t 301ppw@$      sq ~��~-0q ~ q ~�t 302ppw@$      sq ~��~-3�q ~ q ~�t 303ppw@$      sq ~��~-7�q ~ q ~�t 304ppw@$      sq ~��~-;Iq ~ q ~�t 305ppw@$      sq ~��~-?
q ~ q ~�t 306ppw@$      sq ~��~-B�q ~ q ~�t 307ppw@$      sq ~��~-F�q ~ q ~�t 308ppw@$      sq ~��~-JMq ~ q ~�t 309ppw@$      sq ~��{_گq ~ q ~�t 31ppw@$��i�L�sq ~��~-��q ~ q ~�t 310ppw@$      sq ~��~-��q ~ q ~�t 311ppw@$      sq ~��~-�eq ~ q ~�t 312ppw@$      sq ~��~-�&q ~ q ~�t 313ppw@#�i����sq ~��~-��q ~ q ~�t 314ppw@$      sq ~��~-��q ~ q ~�t 315ppw@$      sq ~��~-�iq ~ q ~�t 316ppw@$      sq ~��~-�*q ~ q ~�t 317ppw@$      sq ~��~-��q ~ q ~�t 318ppw@$      sq ~��~-��q ~ q ~�t 319ppw@"J�^�Ysq ~��{_�pq ~ q ~�t 32ppw@$      sq ~��~.Bq ~ q ~�t 320ppw@$      sq ~��~.q ~ q ~�t 321ppw@$      sq ~��~.�q ~ q ~�t 322ppw@$      sq ~��~.�q ~ q ~�t 323ppw@$      sq ~��~. Fq ~ q ~�t 324ppw@$      sq ~��~.$q ~ q ~�t 325ppw@$      sq ~��~.'�q ~ q ~�t 326ppw@$      sq ~��~.+�q ~ q ~�t 327ppw@$      sq ~��~./Jq ~ q ~�t 328ppw@$      sq ~��~.3q ~ q ~�t 329ppw@$      sq ~��{_�1q ~ q ~�t 33ppw@$      sq ~��~.��q ~ q ~�t 330ppw@$      sq ~��~.�bq ~ q ~�t 331ppw@$      sq ~��~.�#q ~ q ~�t 332ppw@$      sq ~��~.��q ~ q ~�t 333ppw@$      sq ~��~.��q ~ q ~�t 334ppw@$      sq ~��~.�fq ~ q ~�t 335ppw@$      sq ~��~.�'q ~ q ~�t 336ppw@$      sq ~��~.��q ~ q ~�t 337ppw@$      sq ~��~.��q ~ q ~�t 338ppw@$      sq ~��~.�jq ~ q ~�t 339ppw@$      sq ~��{_��q ~ q ~�t 34ppw@$`u*D sq ~��~.� q ~ q ~�t 340ppw@$      sq ~��~.��q ~ q ~�t 341ppw@$      sq ~��~/�q ~ q ~�t 342ppw@$      sq ~��~/Cq ~ q ~�t 343ppw@$      sq ~��~/	q ~ q ~�t 344ppw@$      sq ~��~/�q ~ q ~�t 345ppw@$      sq ~��~/�q ~ q ~�t 346ppw@$      sq ~��~/Gq ~ q ~�t 347ppw@$      sq ~��~/q ~ q ~�t 348ppw@$      sq ~��~/�q ~ q ~�t 349ppw@$      sq ~��{_�q ~ q ~�t 35ppw@%�0�g�psq ~��~/n_q ~ q ~�t 350ppw@$      sq ~��~/r q ~ q ~�t 351ppw@$      sq ~��~/u�q ~ q ~�t 352ppw@$      sq ~��~/y�q ~ q ~�t 353ppw@$      sq ~��~/}cq ~ q ~�t 354ppw@$      sq ~��~/�$q ~ q ~�t 355ppw@$      sq ~��~/��q ~ q ~�t 356ppw@$      sq ~��~/��q ~ q ~�t 357ppw@$      sq ~��~/�gq ~ q ~�t 358ppw@$      sq ~��~/�(q ~ q ~�t 359ppw@$      sq ~��{_�tq ~ q ~�t 36ppw@�:NBsq ~��~/�q ~ q ~�t 360ppw@$      sq ~��~/�q ~ q ~�t 361ppw@$      sq ~��~/�@q ~ q ~�t 362ppw@$      sq ~��~/�q ~ q ~�t 363ppw@$      sq ~��~/��q ~ q ~�t 364ppw@$      sq ~��~/��q ~ q ~�t 365ppw@$      sq ~��~/�Dq ~ q ~�t 366ppw@$      sq ~��~/�q ~ q ~�t 367ppw@$      sq ~��~0 �q ~ q ~�t 368ppw@$      sq ~��~0�q ~ q ~�t 369ppw@$      sq ~��{_�5q ~ q ~�t 37ppw@$      sq ~��~0Wq ~ q ~�t 370ppw@$      sq ~��~0Z�q ~ q ~�t 371ppw@$      sq ~��~0^�q ~ q ~�t 372ppw@$      sq ~��~0b`q ~ q ~�t 373ppw@$      sq ~��~0f!q ~ q ~�t 374ppw@$      sq ~��~0i�q ~ q ~�t 375ppw@$      sq ~��~0m�q ~ q ~�t 376ppw@$      sq ~��~0qdq ~ q ~�t 377ppw@$F�\#=�sq ~��~0u%q ~ q ~�t 378ppw@$      sq ~��~0x�q ~ q ~�t 379ppw@$      sq ~��{_��q ~ q ~�t 38ppw@$      sq ~��~0�|q ~ q ~�t 380ppw@$      sq ~��~0�=q ~ q ~�t 381ppw@$      sq ~��~0��q ~ q ~�t 382ppw@$      sq ~��~0ֿq ~ q ~�t 383ppw@$      sq ~��~0ڀq ~ q ~�t 384ppw@$      sq ~��~0�Aq ~ q ~�t 385ppw@$      sq ~��~0�q ~ q ~�t 386ppw@$      sq ~��~0��q ~ q ~�t 387ppw@$      sq ~��~0�q ~ q ~�t 388ppw@$      sq ~��~0�Eq ~ q ~�t 389ppw@$      sq ~��{_��q ~ q ~�t 39ppw@$      sq ~��~1?�q ~ q ~�t 390ppw@$��ɶ�sq ~��~1C�q ~ q ~�t 391ppw@$      sq ~��~1G]q ~ q ~�t 392ppw@$      sq ~��~1Kq ~ q ~�t 393ppw@$      sq ~��~1N�q ~ q ~�t 394ppw@$      sq ~��~1R�q ~ q ~�t 395ppw@$      sq ~��~1Vaq ~ q ~�t 396ppw@$      sq ~��~1Z"q ~ q ~�t 397ppw@$      sq ~��~1]�q ~ q ~�t 398ppw@$      sq ~��~1a�q ~ q ~�t 399ppw@$      sq ~��{H�q ~ q ~�t 4ppw@/g��(�>sq ~��{`KMq ~ q ~�t 40ppw@)�ԋ��sq ~��~;@q ~ q ~�t 400ppw@$      sq ~��~;C�q ~ q ~�t 401ppw@$*a-�Jsq ~��~;G�q ~ q ~�t 402ppw@$      sq ~��~;KHq ~ q ~�t 403ppw@$      sq ~��~;O	q ~ q ~�t 404ppw@$      sq ~��~;R�q ~ q ~�t 405ppw@$      sq ~��~;V�q ~ q ~�t 406ppw@$      sq ~��~;ZLq ~ q ~�t 407ppw@$      sq ~��~;^q ~ q ~�t 408ppw@$      sq ~��~;a�q ~ q ~�t 409ppw@$      sq ~��{`Oq ~ q ~�t 41ppw@)�_��zsq ~��~;�dq ~ q ~�t 410ppw@$      sq ~��~;�%q ~ q ~�t 411ppw@$      sq ~��~;��q ~ q ~�t 412ppw@$      sq ~��~;��q ~ q ~�t 413ppw@$      sq ~��~;�hq ~ q ~�t 414ppw@$      sq ~��~;�)q ~ q ~�t 415ppw@$      sq ~��~;��q ~ q ~�t 416ppw@$      sq ~��~;Ϋq ~ q ~�t 417ppw@$      sq ~��~;�lq ~ q ~�t 418ppw@$      sq ~��~;�-q ~ q ~�t 419ppw@$      sq ~��{`R�q ~ q ~�t 42ppw@'3i���sq ~��~<(�q ~ q ~�t 420ppw@$      sq ~��~<,�q ~ q ~�t 421ppw@%�k԰�sq ~��~<0Eq ~ q ~�t 422ppw@$      sq ~��~<4q ~ q ~�t 423ppw@$      sq ~��~<7�q ~ q ~�t 424ppw@$      sq ~��~<;�q ~ q ~�t 425ppw@%���}B�sq ~��~<?Iq ~ q ~�t 426ppw@$      sq ~��~<C
q ~ q ~�t 427ppw@$      sq ~��~<F�q ~ q ~�t 428ppw@$      sq ~��~<J�q ~ q ~�t 429ppw@$      sq ~��{`V�q ~ q ~�t 43ppw@8��̰�lsq ~��~<�"q ~ q ~�t 430ppw@$      sq ~��~<��q ~ q ~�t 431ppw@$      sq ~��~<��q ~ q ~�t 432ppw@$      sq ~��~<�eq ~ q ~�t 433ppw@$      sq ~��~<�&q ~ q ~�t 434ppw@$      sq ~��~<��q ~ q ~�t 435ppw@$      sq ~��~<��q ~ q ~�t 436ppw@$      sq ~��~<�iq ~ q ~�t 437ppw@$      sq ~��~<�*q ~ q ~�t 438ppw@$      sq ~��~<��q ~ q ~�t 439ppw@$      sq ~��{`ZQq ~ q ~�t 44ppw@$      sq ~��~=�q ~ q ~�t 440ppw@$      sq ~��~=Bq ~ q ~�t 441ppw@$      sq ~��~=q ~ q ~�t 442ppw@$      sq ~��~=�q ~ q ~�t 443ppw@$      sq ~��~= �q ~ q ~�t 444ppw@$      sq ~��~=$Fq ~ q ~�t 445ppw@$      sq ~��~=(q ~ q ~�t 446ppw@$      sq ~��~=+�q ~ q ~�t 447ppw@$      sq ~��~=/�q ~ q ~�t 448ppw@$      sq ~��~=3Jq ~ q ~�t 449ppw@#3^-��sq ~��{`^q ~ q ~�t 45ppw@&φ
6�sq ~��~=��q ~ q ~�t 450ppw@$      sq ~��~=��q ~ q ~�t 451ppw@$      sq ~��~=�bq ~ q ~�t 452ppw@$      sq ~��~=�#q ~ q ~�t 453ppw@$      sq ~��~=��q ~ q ~�t 454ppw@$      sq ~��~=��q ~ q ~�t 455ppw@$      sq ~��~=�fq ~ q ~�t 456ppw@"5w��sq ~��~=�'q ~ q ~�t 457ppw@$      sq ~��~=��q ~ q ~�t 458ppw@$      sq ~��~=��q ~ q ~�t 459ppw@$      sq ~��{`a�q ~ q ~�t 46ppw@&�Idc�sq ~��~=�?q ~ q ~�t 460ppw@$      sq ~��~=� q ~ q ~�t 461ppw@$      sq ~��~>�q ~ q ~�t 462ppw@$      sq ~��~>�q ~ q ~�t 463ppw@$      sq ~��~>	Cq ~ q ~�t 464ppw@$      sq ~��~>q ~ q ~�t 465ppw@$      sq ~��~>�q ~ q ~�t 466ppw@$      sq ~��~>�q ~ q ~�t 467ppw@$      sq ~��~>Gq ~ q ~�t 468ppw@$      sq ~��~>q ~ q ~�t 469ppw@$      sq ~��{`e�q ~ q ~�t 47ppw@"�}/��sq ~��~>n�q ~ q ~�t 470ppw@$      sq ~��~>r_q ~ q ~�t 471ppw@$      sq ~��~>v q ~ q ~�t 472ppw@$      sq ~��~>y�q ~ q ~�t 473ppw@$      sq ~��~>}�q ~ q ~�t 474ppw@$      sq ~��~>�cq ~ q ~�t 475ppw@$      sq ~��~>�$q ~ q ~�t 476ppw@$      sq ~��~>��q ~ q ~�t 477ppw@$      sq ~��~>��q ~ q ~�t 478ppw@$      sq ~��~>�gq ~ q ~�t 479ppw@$      sq ~��{`iUq ~ q ~�t 48ppw@)*��sq ~��~>��q ~ q ~�t 480ppw@$      sq ~��~>�q ~ q ~�t 481ppw@$      sq ~��~>�q ~ q ~�t 482ppw@$      sq ~��~>�@q ~ q ~�t 483ppw@$      sq ~��~>�q ~ q ~�t 484ppw@$      sq ~��~>��q ~ q ~�t 485ppw@$      sq ~��~>��q ~ q ~�t 486ppw@$      sq ~��~>�Dq ~ q ~�t 487ppw@$      sq ~��~?q ~ q ~�t 488ppw@$      sq ~��~?�q ~ q ~�t 489ppw@$      sq ~��{`mq ~ q ~�t 49ppw@&��+Asq ~��~?W\q ~ q ~�t 490ppw@#���*�sq ~��~?[q ~ q ~�t 491ppw@$      sq ~��~?^�q ~ q ~�t 492ppw@$      sq ~��~?b�q ~ q ~�t 493ppw@$      sq ~��~?f`q ~ q ~�t 494ppw@$      sq ~��~?j!q ~ q ~�t 495ppw@$      sq ~��~?m�q ~ q ~�t 496ppw@$      sq ~��~?q�q ~ q ~�t 497ppw@$      sq ~��~?udq ~ q ~�t 498ppw@$      sq ~��~?y%q ~ q ~�t 499ppw@$      sq ~��{H��q ~ q ~�t 5ppw@&����]2sq ~��{`��q ~ q ~�t 50ppw@~Xl�uCsq ~��~IW�q ~ q ~�t 500ppw@$      sq ~��~I[Gq ~ q ~�t 501ppw@$      sq ~��~I_q ~ q ~�t 502ppw@$      sq ~��~Ib�q ~ q ~�t 503ppw@$      sq ~��~If�q ~ q ~�t 504ppw@$      sq ~��~IjKq ~ q ~�t 505ppw@$      sq ~��~Inq ~ q ~�t 506ppw@$      sq ~��~Iq�q ~ q ~�t 507ppw@$      sq ~��~Iu�q ~ q ~�t 508ppw@$      sq ~��~IyOq ~ q ~�t 509ppw@$      sq ~��{`�mq ~ q ~�t 51ppw@0��RZY�sq ~��~I��q ~ q ~�t 510ppw@$      sq ~��~IϦq ~ q ~�t 511ppw@$      sq ~��~I�gq ~ q ~�t 512ppw@$      sq ~��~I�(q ~ q ~�t 513ppw@$      sq ~��~I��q ~ q ~�t 514ppw@$      sq ~��~Iުq ~ q ~�t 515ppw@$      sq ~��~I�kq ~ q ~�t 516ppw@$      sq ~��~I�,q ~ q ~�t 517ppw@$      sq ~��~I��q ~ q ~�t 518ppw@$      sq ~��~I�q ~ q ~�t 519ppw@$      sq ~��{`�.q ~ q ~�t 52ppw@$      sq ~��~J@Dq ~ q ~�t 520ppw@$      sq ~��~JDq ~ q ~�t 521ppw@$      sq ~��~JG�q ~ q ~�t 522ppw@$      sq ~��~JK�q ~ q ~�t 523ppw@$      sq ~��~JOHq ~ q ~�t 524ppw@$&L��@sq ~��~JS	q ~ q ~�t 525ppw@$      sq ~��~JV�q ~ q ~�t 526ppw@$      sq ~��~JZ�q ~ q ~�t 527ppw@$      sq ~��~J^Lq ~ q ~�t 528ppw@$      sq ~��~Jbq ~ q ~�t 529ppw@$      sq ~��{`��q ~ q ~�t 53ppw@#>��sq ~��~J��q ~ q ~�t 530ppw@$      sq ~��~J�dq ~ q ~�t 531ppw@$      sq ~��~J�%q ~ q ~�t 532ppw@$      sq ~��~J��q ~ q ~�t 533ppw@$      sq ~��~Jçq ~ q ~�t 534ppw@$      sq ~��~J�hq ~ q ~�t 535ppw@$      sq ~��~J�)q ~ q ~�t 536ppw@$      sq ~��~J��q ~ q ~�t 537ppw@$      sq ~��~Jҫq ~ q ~�t 538ppw@$      sq ~��~J�lq ~ q ~�t 539ppw@$      sq ~��{`ΰq ~ q ~�t 54ppw@$      sq ~��~K)q ~ q ~�t 540ppw@$      sq ~��~K,�q ~ q ~�t 541ppw@$      sq ~��~K0�q ~ q ~�t 542ppw@$      sq ~��~K4Eq ~ q ~�t 543ppw@$      sq ~��~K8q ~ q ~�t 544ppw@$      sq ~��~K;�q ~ q ~�t 545ppw@$      sq ~��~K?�q ~ q ~�t 546ppw@$      sq ~��~KCIq ~ q ~�t 547ppw@$      sq ~��~KG
q ~ q ~�t 548ppw@$      sq ~��~KJ�q ~ q ~�t 549ppw@$      sq ~��{`�qq ~ q ~�t 55ppw@$      sq ~��~K�aq ~ q ~�t 550ppw@$      sq ~��~K�"q ~ q ~�t 551ppw@$      sq ~��~K��q ~ q ~�t 552ppw@$      sq ~��~K��q ~ q ~�t 553ppw@$      sq ~��~K�eq ~ q ~�t 554ppw@$      sq ~��~K�&q ~ q ~�t 555ppw@$      sq ~��~K��q ~ q ~�t 556ppw@$      sq ~��~K��q ~ q ~�t 557ppw@$      sq ~��~K�iq ~ q ~�t 558ppw@$      sq ~��~K�*q ~ q ~�t 559ppw@$      sq ~��{`�2q ~ q ~�t 56ppw@#�2�?sq ~��~L�q ~ q ~�t 560ppw@$      sq ~��~L�q ~ q ~�t 561ppw@$      sq ~��~LBq ~ q ~�t 562ppw@$      sq ~��~Lq ~ q ~�t 563ppw@$      sq ~��~L �q ~ q ~�t 564ppw@$      sq ~��~L$�q ~ q ~�t 565ppw@$      sq ~��~L(Fq ~ q ~�t 566ppw@$      sq ~��~L,q ~ q ~�t 567ppw@$      sq ~��~L/�q ~ q ~�t 568ppw@$      sq ~��~L3�q ~ q ~�t 569ppw@$      sq ~��{`��q ~ q ~�t 57ppw@$      sq ~��~L�q ~ q ~�t 570ppw@$      sq ~��~L��q ~ q ~�t 571ppw@$      sq ~��~L��q ~ q ~�t 572ppw@$      sq ~��~L�bq ~ q ~�t 573ppw@$      sq ~��~L�#q ~ q ~�t 574ppw@$      sq ~��~L��q ~ q ~�t 575ppw@$      sq ~��~L��q ~ q ~�t 576ppw@$      sq ~��~L�fq ~ q ~�t 577ppw@$      sq ~��~L�'q ~ q ~�t 578ppw@$      sq ~��~L��q ~ q ~�t 579ppw@$      sq ~��{`ݴq ~ q ~�t 58ppw@6C����sq ~��~L�~q ~ q ~�t 580ppw@$      sq ~��~L�?q ~ q ~�t 581ppw@$      sq ~��~M q ~ q ~�t 582ppw@$      sq ~��~M�q ~ q ~�t 583ppw@$      sq ~��~M	�q ~ q ~�t 584ppw@$      sq ~��~MCq ~ q ~�t 585ppw@$      sq ~��~Mq ~ q ~�t 586ppw@$      sq ~��~M�q ~ q ~�t 587ppw@$      sq ~��~M�q ~ q ~�t 588ppw@$      sq ~��~MGq ~ q ~�t 589ppw@$      sq ~��{`�uq ~ q ~�t 59ppw@&a���O�sq ~��~Mn�q ~ q ~�t 590ppw@$      sq ~��~Mr�q ~ q ~�t 591ppw@$      sq ~��~Mv_q ~ q ~�t 592ppw@$      sq ~��~Mz q ~ q ~�t 593ppw@$      sq ~��~M}�q ~ q ~�t 594ppw@$      sq ~��~M��q ~ q ~�t 595ppw@$      sq ~��~M�cq ~ q ~�t 596ppw@$      sq ~��~M�$q ~ q ~�t 597ppw@$      sq ~��~M��q ~ q ~�t 598ppw@$      sq ~��~M��q ~ q ~�t 599ppw@$      sq ~��{H��q ~ q ~�t 6ppw@?iݝ��sq ~��{a4q ~ q ~�t 60ppw@$      sq ~��~Woq ~ q ~�t 600ppw@$      sq ~��~Wr�q ~ q ~�t 601ppw@$      sq ~��~Wv�q ~ q ~�t 602ppw@$      sq ~��~WzJq ~ q ~�t 603ppw@$      sq ~��~W~q ~ q ~�t 604ppw@$      sq ~��~W��q ~ q ~�t 605ppw@$      sq ~��~W��q ~ q ~�t 606ppw@$      sq ~��~W�Nq ~ q ~�t 607ppw@$      sq ~��~W�q ~ q ~�t 608ppw@$      sq ~��~W��q ~ q ~�t 609ppw@$      sq ~��{a7�q ~ q ~�t 61ppw@&V6��sq ~��~W�fq ~ q ~�t 610ppw@$      sq ~��~W�'q ~ q ~�t 611ppw@$      sq ~��~W��q ~ q ~�t 612ppw@$      sq ~��~W�q ~ q ~�t 613ppw@$      sq ~��~W�jq ~ q ~�t 614ppw@$      sq ~��~W�+q ~ q ~�t 615ppw@$      sq ~��~W��q ~ q ~�t 616ppw@$      sq ~��~W��q ~ q ~�t 617ppw@$      sq ~��~Xnq ~ q ~�t 618ppw@$      sq ~��~X/q ~ q ~�t 619ppw@$      sq ~��{a;�q ~ q ~�t 62ppw@$*�$F�Nsq ~��~XW�q ~ q ~�t 620ppw@$      sq ~��~X[�q ~ q ~�t 621ppw@$      sq ~��~X_Gq ~ q ~�t 622ppw@$      sq ~��~Xcq ~ q ~�t 623ppw@$      sq ~��~Xf�q ~ q ~�t 624ppw@$      sq ~��~Xj�q ~ q ~�t 625ppw@$      sq ~��~XnKq ~ q ~�t 626ppw@$      sq ~��~Xrq ~ q ~�t 627ppw@$      sq ~��~Xu�q ~ q ~�t 628ppw@$      sq ~��~Xy�q ~ q ~�t 629ppw@$      sq ~��{a?Nq ~ q ~�t 63ppw@&�'w�sq ~��~X�$q ~ q ~�t 630ppw@$      sq ~��~X��q ~ q ~�t 631ppw@$      sq ~��~XӦq ~ q ~�t 632ppw@$      sq ~��~X�gq ~ q ~�t 633ppw@$      sq ~��~X�(q ~ q ~�t 634ppw@$      sq ~��~X��q ~ q ~�t 635ppw@$      sq ~��~X�q ~ q ~�t 636ppw@$      sq ~��~X�kq ~ q ~�t 637ppw@$      sq ~��~X�,q ~ q ~�t 638ppw@$      sq ~��~X��q ~ q ~�t 639ppw@$      sq ~��{aCq ~ q ~�t 64ppw@$      sq ~��~Y@�q ~ q ~�t 640ppw@$      sq ~��~YDDq ~ q ~�t 641ppw@$      sq ~��~YHq ~ q ~�t 642ppw@$      sq ~��~YK�q ~ q ~�t 643ppw@$      sq ~��~YO�q ~ q ~�t 644ppw@$      sq ~��~YSHq ~ q ~�t 645ppw@$      sq ~��~YW	q ~ q ~�t 646ppw@$      sq ~��~YZ�q ~ q ~�t 647ppw@$      sq ~��~Y^�q ~ q ~�t 648ppw@$      sq ~��~YbLq ~ q ~�t 649ppw@$      sq ~��{aF�q ~ q ~�t 65ppw@0v�Ok��sq ~��~Y��q ~ q ~�t 650ppw@$      sq ~��~Y��q ~ q ~�t 651ppw@$      sq ~��~Y�dq ~ q ~�t 652ppw@$      sq ~��~Y�%q ~ q ~�t 653ppw@$      sq ~��~Y��q ~ q ~�t 654ppw@$      sq ~��~Yǧq ~ q ~�t 655ppw@$      sq ~��~Y�hq ~ q ~�t 656ppw@$      sq ~��~Y�)q ~ q ~�t 657ppw@$      sq ~��~Y��q ~ q ~�t 658ppw@$      sq ~��~Y֫q ~ q ~�t 659ppw@$      sq ~��{aJ�q ~ q ~�t 66ppw@$      sq ~��~Z)Aq ~ q ~�t 660ppw@$      sq ~��~Z-q ~ q ~�t 661ppw@$      sq ~��~Z0�q ~ q ~�t 662ppw@$      sq ~��~Z4�q ~ q ~�t 663ppw@$      sq ~��~Z8Eq ~ q ~�t 664ppw@$      sq ~��~Z<q ~ q ~�t 665ppw@$      sq ~��~Z?�q ~ q ~�t 666ppw@$      sq ~��~ZC�q ~ q ~�t 667ppw@$      sq ~��~ZGIq ~ q ~�t 668ppw@$      sq ~��~ZK
q ~ q ~�t 669ppw@$      sq ~��{aNRq ~ q ~�t 67ppw@%��P	�sq ~��~Z��q ~ q ~�t 670ppw@$      sq ~��~Z�aq ~ q ~�t 671ppw@$      sq ~��~Z�"q ~ q ~�t 672ppw@$      sq ~��~Z��q ~ q ~�t 673ppw@$      sq ~��~Z��q ~ q ~�t 674ppw@$      sq ~��~Z�eq ~ q ~�t 675ppw@$      sq ~��~Z�&q ~ q ~�t 676ppw@$      sq ~��~Z��q ~ q ~�t 677ppw@$      sq ~��~Z��q ~ q ~�t 678ppw@$      sq ~��~Z�iq ~ q ~�t 679ppw@$      sq ~��{aRq ~ q ~�t 68ppw@/v8p�}�sq ~��~[�q ~ q ~�t 680ppw@$      sq ~��~[�q ~ q ~�t 681ppw@$      sq ~��~[�q ~ q ~�t 682ppw@$      sq ~��~[Bq ~ q ~�t 683ppw@$      sq ~��~[!q ~ q ~�t 684ppw@$      sq ~��~[$�q ~ q ~�t 685ppw@$      sq ~��~[(�q ~ q ~�t 686ppw@$      sq ~��~[,Fq ~ q ~�t 687ppw@#�l��sq ~��~[0q ~ q ~�t 688ppw@$      sq ~��~[3�q ~ q ~�t 689ppw@$      sq ~��{aU�q ~ q ~�t 69ppw@ _eq�sq ~��~[�^q ~ q ~�t 690ppw@$      sq ~��~[�q ~ q ~�t 691ppw@$      sq ~��~[��q ~ q ~�t 692ppw@$      sq ~��~[��q ~ q ~�t 693ppw@$      sq ~��~[�bq ~ q ~�t 694ppw@$      sq ~��~[�#q ~ q ~�t 695ppw@$      sq ~��~[��q ~ q ~�t 696ppw@$      sq ~��~[��q ~ q ~�t 697ppw@$      sq ~��~[�fq ~ q ~�t 698ppw@$      sq ~��~[�'q ~ q ~�t 699ppw@$      sq ~��{H�Hq ~ q ~�t 7ppw@'�37�sq ~��{a�jq ~ q ~�t 70ppw@$      sq ~��~e��q ~ q ~�t 700ppw@$      sq ~��~e�Iq ~ q ~�t 701ppw@$      sq ~��~e�
q ~ q ~�t 702ppw@$      sq ~��~e��q ~ q ~�t 703ppw@$      sq ~��~e��q ~ q ~�t 704ppw@$      sq ~��~e�Mq ~ q ~�t 705ppw@$      sq ~��~e�q ~ q ~�t 706ppw@$      sq ~��~e��q ~ q ~�t 707ppw@$      sq ~��~e��q ~ q ~�t 708ppw@$      sq ~��~e�Qq ~ q ~�t 709ppw@$      sq ~��{a�+q ~ q ~�t 71ppw@$      sq ~��~e��q ~ q ~�t 710ppw@$      sq ~��~e��q ~ q ~�t 711ppw@$      sq ~��~fiq ~ q ~�t 712ppw@$      sq ~��~f*q ~ q ~�t 713ppw@$      sq ~��~f	�q ~ q ~�t 714ppw@$      sq ~��~f�q ~ q ~�t 715ppw@$      sq ~��~fmq ~ q ~�t 716ppw@$      sq ~��~f.q ~ q ~�t 717ppw@$      sq ~��~f�q ~ q ~�t 718ppw@$      sq ~��~f�q ~ q ~�t 719ppw@$      sq ~��{a��q ~ q ~�t 72ppw@$      sq ~��~foFq ~ q ~�t 720ppw@$      sq ~��~fsq ~ q ~�t 721ppw@$      sq ~��~fv�q ~ q ~�t 722ppw@$      sq ~��~fz�q ~ q ~�t 723ppw@$      sq ~��~f~Jq ~ q ~�t 724ppw@$      sq ~��~f�q ~ q ~�t 725ppw@$      sq ~��~f��q ~ q ~�t 726ppw@$      sq ~��~f��q ~ q ~�t 727ppw@$      sq ~��~f�Nq ~ q ~�t 728ppw@$      sq ~��~f�q ~ q ~�t 729ppw@$      sq ~��{a��q ~ q ~�t 73ppw@$      sq ~��~f�q ~ q ~�t 730ppw@$      sq ~��~f�fq ~ q ~�t 731ppw@$      sq ~��~f�'q ~ q ~�t 732ppw@$      sq ~��~f��q ~ q ~�t 733ppw@$      sq ~��~f�q ~ q ~�t 734ppw@$      sq ~��~f�jq ~ q ~�t 735ppw@$      sq ~��~f�+q ~ q ~�t 736ppw@#��Ё�sq ~��~f��q ~ q ~�t 737ppw@$      sq ~��~g�q ~ q ~�t 738ppw@$      sq ~��~gnq ~ q ~�t 739ppw@#ٳ�:�sq ~��{a�nq ~ q ~�t 74ppw@�����msq ~��~gXq ~ q ~�t 740ppw@$      sq ~��~g[�q ~ q ~�t 741ppw@$      sq ~��~g_�q ~ q ~�t 742ppw@$      sq ~��~gcGq ~ q ~�t 743ppw@$      sq ~��~ggq ~ q ~�t 744ppw@$      sq ~��~gj�q ~ q ~�t 745ppw@$      sq ~��~gn�q ~ q ~�t 746ppw@$      sq ~��~grKq ~ q ~�t 747ppw@$      sq ~��~gvq ~ q ~�t 748ppw@$      sq ~��~gy�q ~ q ~�t 749ppw@$      sq ~��{a�/q ~ q ~�t 75ppw@)ꑷ(�lsq ~��~g�cq ~ q ~�t 750ppw@$      sq ~��~g�$q ~ q ~�t 751ppw@$      sq ~��~g��q ~ q ~�t 752ppw@$      sq ~��~gצq ~ q ~�t 753ppw@$      sq ~��~g�gq ~ q ~�t 754ppw@$      sq ~��~g�(q ~ q ~�t 755ppw@$      sq ~��~g��q ~ q ~�t 756ppw@$      sq ~��~g�q ~ q ~�t 757ppw@$      sq ~��~g�kq ~ q ~�t 758ppw@$      sq ~��~g�,q ~ q ~�t 759ppw@$      sq ~��{a��q ~ q ~�t 76ppw@$      sq ~��~h@�q ~ q ~�t 760ppw@$      sq ~��~hD�q ~ q ~�t 761ppw@$      sq ~��~hHDq ~ q ~�t 762ppw@$      sq ~��~hLq ~ q ~�t 763ppw@$      sq ~��~hO�q ~ q ~�t 764ppw@$      sq ~��~hS�q ~ q ~�t 765ppw@$      sq ~��~hWHq ~ q ~�t 766ppw@$      sq ~��~h[	q ~ q ~�t 767ppw@$      sq ~��~h^�q ~ q ~�t 768ppw@$      sq ~��~hb�q ~ q ~�t 769ppw@$      sq ~��{a±q ~ q ~�t 77ppw@"��d`�sq ~��~h�!q ~ q ~�t 770ppw@$      sq ~��~h��q ~ q ~�t 771ppw@$      sq ~��~h��q ~ q ~�t 772ppw@$      sq ~��~h�dq ~ q ~�t 773ppw@$      sq ~��~h�%q ~ q ~�t 774ppw@$      sq ~��~h��q ~ q ~�t 775ppw@$      sq ~��~h˧q ~ q ~�t 776ppw@$      sq ~��~h�hq ~ q ~�t 777ppw@$      sq ~��~h�)q ~ q ~�t 778ppw@$      sq ~��~h��q ~ q ~�t 779ppw@$      sq ~��{a�rq ~ q ~�t 78ppw@$      sq ~��~i)�q ~ q ~�t 780ppw@$      sq ~��~i-Aq ~ q ~�t 781ppw@$      sq ~��~i1q ~ q ~�t 782ppw@$      sq ~��~i4�q ~ q ~�t 783ppw@$      sq ~��~i8�q ~ q ~�t 784ppw@$      sq ~��~i<Eq ~ q ~�t 785ppw@$      sq ~��~i@q ~ q ~�t 786ppw@$      sq ~��~iC�q ~ q ~�t 787ppw@$      sq ~��~iG�q ~ q ~�t 788ppw@$      sq ~��~iKIq ~ q ~�t 789ppw@$      sq ~��{a�3q ~ q ~�t 79ppw@#�^e�R�sq ~��~i��q ~ q ~�t 790ppw@$      sq ~��~i��q ~ q ~�t 791ppw@$      sq ~��~i�aq ~ q ~�t 792ppw@$      sq ~��~i�"q ~ q ~�t 793ppw@$      sq ~��~i��q ~ q ~�t 794ppw@$      sq ~��~i��q ~ q ~�t 795ppw@$      sq ~��~i�eq ~ q ~�t 796ppw@$      sq ~��~i�&q ~ q ~�t 797ppw@$      sq ~��~i��q ~ q ~�t 798ppw@$      sq ~��~i��q ~ q ~�t 799ppw@$      sq ~��{H�	q ~ q ~�t 8ppw@$      sq ~��{b�q ~ q ~�t 80ppw@$      sq ~��~s�	q ~ q ~�t 800ppw@$      sq ~��~s��q ~ q ~�t 801ppw@$      sq ~��~s��q ~ q ~�t 802ppw@$      sq ~��~s�Lq ~ q ~�t 803ppw@$>�(R=�sq ~��~s�q ~ q ~�t 804ppw@$      sq ~��~s��q ~ q ~�t 805ppw@$      sq ~��~s��q ~ q ~�t 806ppw@$      sq ~��~s�Pq ~ q ~�t 807ppw@$      sq ~��~s�q ~ q ~�t 808ppw@$      sq ~��~s��q ~ q ~�t 809ppw@$      sq ~��{b �q ~ q ~�t 81ppw@$      sq ~��~thq ~ q ~�t 810ppw@$      sq ~��~t)q ~ q ~�t 811ppw@$      sq ~��~t�q ~ q ~�t 812ppw@$      sq ~��~t�q ~ q ~�t 813ppw@$      sq ~��~t!lq ~ q ~�t 814ppw@$      sq ~��~t%-q ~ q ~�t 815ppw@$��BB�sq ~��~t(�q ~ q ~�t 816ppw@$      sq ~��~t,�q ~ q ~�t 817ppw@$      sq ~��~t0pq ~ q ~�t 818ppw@$      sq ~��~t41q ~ q ~�t 819ppw@$      sq ~��{b$Kq ~ q ~�t 82ppw@$      sq ~��~t��q ~ q ~�t 820ppw@$      sq ~��~t��q ~ q ~�t 821ppw@$      sq ~��~t�Iq ~ q ~�t 822ppw@$      sq ~��~t�
q ~ q ~�t 823ppw@$      sq ~��~t��q ~ q ~�t 824ppw@$      sq ~��~t��q ~ q ~�t 825ppw@$      sq ~��~t�Mq ~ q ~�t 826ppw@$      sq ~��~t�q ~ q ~�t 827ppw@$      sq ~��~t��q ~ q ~�t 828ppw@$      sq ~��~t��q ~ q ~�t 829ppw@$      sq ~��{b(q ~ q ~�t 83ppw@�D���sq ~��~t�&q ~ q ~�t 830ppw@&����%Bsq ~��~t��q ~ q ~�t 831ppw@$      sq ~��~u�q ~ q ~�t 832ppw@$      sq ~��~uiq ~ q ~�t 833ppw@$      sq ~��~u
*q ~ q ~�t 834ppw@$      sq ~��~u�q ~ q ~�t 835ppw@$      sq ~��~u�q ~ q ~�t 836ppw@$      sq ~��~umq ~ q ~�t 837ppw@$      sq ~��~u.q ~ q ~�t 838ppw@$      sq ~��~u�q ~ q ~�t 839ppw@$      sq ~��{b+�q ~ q ~�t 84ppw@$e{i�sq ~��~uo�q ~ q ~�t 840ppw@$      sq ~��~usFq ~ q ~�t 841ppw@$      sq ~��~uwq ~ q ~�t 842ppw@$      sq ~��~uz�q ~ q ~�t 843ppw@$      sq ~��~u~�q ~ q ~�t 844ppw@$      sq ~��~u�Jq ~ q ~�t 845ppw@$      sq ~��~u�q ~ q ~�t 846ppw@$      sq ~��~u��q ~ q ~�t 847ppw@$      sq ~��~u��q ~ q ~�t 848ppw@$      sq ~��~u�Nq ~ q ~�t 849ppw@$      sq ~��{b/�q ~ q ~�t 85ppw@$      sq ~��~u��q ~ q ~�t 850ppw@$      sq ~��~u�q ~ q ~�t 851ppw@"��r
sq ~��~u�fq ~ q ~�t 852ppw@$      sq ~��~u�'q ~ q ~�t 853ppw@$      sq ~��~u��q ~ q ~�t 854ppw@$      sq ~��~u��q ~ q ~�t 855ppw@$      sq ~��~u�jq ~ q ~�t 856ppw@"��a�5sq ~��~u�+q ~ q ~�t 857ppw@$      sq ~��~v�q ~ q ~�t 858ppw@$      sq ~��~v�q ~ q ~�t 859ppw@$      sq ~��{b3Oq ~ q ~�t 86ppw@2ڐ��?"sq ~��~vXCq ~ q ~�t 860ppw@$      sq ~��~v\q ~ q ~�t 861ppw@$      sq ~��~v_�q ~ q ~�t 862ppw@$      sq ~��~vc�q ~ q ~�t 863ppw@#�B5_Z�sq ~��~vgGq ~ q ~�t 864ppw@$      sq ~��~vkq ~ q ~�t 865ppw@$      sq ~��~vn�q ~ q ~�t 866ppw@$      sq ~��~vr�q ~ q ~�t 867ppw@$      sq ~��~vvKq ~ q ~�t 868ppw@$      sq ~��~vzq ~ q ~�t 869ppw@$      sq ~��{b7q ~ q ~�t 87ppw@$      sq ~��~v̢q ~ q ~�t 870ppw@$      sq ~��~v�cq ~ q ~�t 871ppw@$      sq ~��~v�$q ~ q ~�t 872ppw@$      sq ~��~v��q ~ q ~�t 873ppw@$      sq ~��~vۦq ~ q ~�t 874ppw@$      sq ~��~v�gq ~ q ~�t 875ppw@$      sq ~��~v�(q ~ q ~�t 876ppw@$      sq ~��~v��q ~ q ~�t 877ppw@$      sq ~��~v�q ~ q ~�t 878ppw@$      sq ~��~v�kq ~ q ~�t 879ppw@$      sq ~��{b:�q ~ q ~�t 88ppw@ ֡r�X�sq ~��~wAq ~ q ~�t 880ppw@$      sq ~��~wD�q ~ q ~�t 881ppw@$      sq ~��~wH�q ~ q ~�t 882ppw@$      sq ~��~wLDq ~ q ~�t 883ppw@$      sq ~��~wPq ~ q ~�t 884ppw@$      sq ~��~wS�q ~ q ~�t 885ppw@$      sq ~��~wW�q ~ q ~�t 886ppw@$      sq ~��~w[Hq ~ q ~�t 887ppw@$      sq ~��~w_	q ~ q ~�t 888ppw@%��<\�sq ~��~wb�q ~ q ~�t 889ppw@$      sq ~��{b>�q ~ q ~�t 89ppw@%��+Lsq ~��~w�`q ~ q ~�t 890ppw@$      sq ~��~w�!q ~ q ~�t 891ppw@$      sq ~��~w��q ~ q ~�t 892ppw@$      sq ~��~w��q ~ q ~�t 893ppw@$      sq ~��~w�dq ~ q ~�t 894ppw@$      sq ~��~w�%q ~ q ~�t 895ppw@$      sq ~��~w��q ~ q ~�t 896ppw@$      sq ~��~wϧq ~ q ~�t 897ppw@$      sq ~��~w�hq ~ q ~�t 898ppw@$      sq ~��~w�)q ~ q ~�t 899ppw@$      sq ~��{H��q ~ q ~�t 9ppw@$      sq ~��{b�(q ~ q ~�t 90ppw@$      sq ~��~���q ~ q ~�t 900ppw@$      sq ~��~��Kq ~ q ~�t 901ppw@$      sq ~��~��q ~ q ~�t 902ppw@$      sq ~��~���q ~ q ~�t 903ppw@$      sq ~��~�Ďq ~ q ~�t 904ppw@$      sq ~��~��Oq ~ q ~�t 905ppw@$      sq ~��~��q ~ q ~�t 906ppw@$      sq ~��~���q ~ q ~�t 907ppw@$      sq ~��~�Ӓq ~ q ~�t 908ppw@$      sq ~��~��Sq ~ q ~�t 909ppw@$      sq ~��{b��q ~ q ~�t 91ppw@)94Go�sq ~��~�)�q ~ q ~�t 910ppw@$      sq ~��~�-�q ~ q ~�t 911ppw@$      sq ~��~�1kq ~ q ~�t 912ppw@$      sq ~��~�5,q ~ q ~�t 913ppw@$      sq ~��~�8�q ~ q ~�t 914ppw@$      sq ~��~�<�q ~ q ~�t 915ppw@$      sq ~��~�@oq ~ q ~�t 916ppw@$      sq ~��~�D0q ~ q ~�t 917ppw@$      sq ~��~�G�q ~ q ~�t 918ppw@$      sq ~��~�K�q ~ q ~�t 919ppw@$      sq ~��{b��q ~ q ~�t 92ppw@��Esq ~��~��Hq ~ q ~�t 920ppw@$      sq ~��~��	q ~ q ~�t 921ppw@$      sq ~��~���q ~ q ~�t 922ppw@$      sq ~��~���q ~ q ~�t 923ppw@$      sq ~��~��Lq ~ q ~�t 924ppw@$      sq ~��~��q ~ q ~�t 925ppw@$      sq ~��~���q ~ q ~�t 926ppw@$      sq ~��~���q ~ q ~�t 927ppw@$      sq ~��~��Pq ~ q ~�t 928ppw@$      sq ~��~��q ~ q ~�t 929ppw@$      sq ~��{b�kq ~ q ~�t 93ppw@&n��:ssq ~��~��q ~ q ~�t 930ppw@$      sq ~��~�hq ~ q ~�t 931ppw@$      sq ~��~�)q ~ q ~�t 932ppw@$      sq ~��~��q ~ q ~�t 933ppw@$      sq ~��~�!�q ~ q ~�t 934ppw@$      sq ~��~�%lq ~ q ~�t 935ppw@$      sq ~��~�)-q ~ q ~�t 936ppw@$      sq ~��~�,�q ~ q ~�t 937ppw@$      sq ~��~�0�q ~ q ~�t 938ppw@$      sq ~��~�4pq ~ q ~�t 939ppw@$      sq ~��{b�,q ~ q ~�t 94ppw@!^ƪT��sq ~��~��q ~ q ~�t 940ppw@$      sq ~��~���q ~ q ~�t 941ppw@$#�a�
sq ~��~���q ~ q ~�t 942ppw@$      sq ~��~��Iq ~ q ~�t 943ppw@$      sq ~��~��
q ~ q ~�t 944ppw@$      sq ~��~���q ~ q ~�t 945ppw@$      sq ~��~���q ~ q ~�t 946ppw@$      sq ~��~��Mq ~ q ~�t 947ppw@$      sq ~��~��q ~ q ~�t 948ppw@$      sq ~��~���q ~ q ~�t 949ppw@$      sq ~��{b��q ~ q ~�t 95ppw?�3�_�sq ~��~��eq ~ q ~�t 950ppw@$      sq ~��~��&q ~ q ~�t 951ppw@$      sq ~��~��q ~ q ~�t 952ppw@$      sq ~��~��q ~ q ~�t 953ppw@$      sq ~��~�
iq ~ q ~�t 954ppw@$      sq ~��~�*q ~ q ~�t 955ppw@$      sq ~��~��q ~ q ~�t 956ppw@$      sq ~��~��q ~ q ~�t 957ppw@$      sq ~��~�mq ~ q ~�t 958ppw@$      sq ~��~�.q ~ q ~�t 959ppw@$      sq ~��{b��q ~ q ~�t 96ppw@$%Cє��sq ~��~�o�q ~ q ~�t 960ppw@$      sq ~��~�s�q ~ q ~�t 961ppw@$      sq ~��~�wFq ~ q ~�t 962ppw@$      sq ~��~�{q ~ q ~�t 963ppw@$      sq ~��~�~�q ~ q ~�t 964ppw@$      sq ~��~���q ~ q ~�t 965ppw@$      sq ~��~��Jq ~ q ~�t 966ppw@$      sq ~��~��q ~ q ~�t 967ppw@$      sq ~��~���q ~ q ~�t 968ppw@$      sq ~��~���q ~ q ~�t 969ppw@$      sq ~��{b�oq ~ q ~�t 97ppw@$      sq ~��~��#q ~ q ~�t 970ppw@$      sq ~��~���q ~ q ~�t 971ppw@$      sq ~��~��q ~ q ~�t 972ppw@$      sq ~��~��fq ~ q ~�t 973ppw@$      sq ~��~��'q ~ q ~�t 974ppw@$      sq ~��~���q ~ q ~�t 975ppw@$      sq ~��~���q ~ q ~�t 976ppw@$      sq ~��~��jq ~ q ~�t 977ppw@$      sq ~��~�+q ~ q ~�t 978ppw@$      sq ~��~��q ~ q ~�t 979ppw@$      sq ~��{b�0q ~ q ~�t 98ppw@.;1�6sq ~��~�X�q ~ q ~�t 980ppw@$      sq ~��~�\Cq ~ q ~�t 981ppw@$      sq ~��~�`q ~ q ~�t 982ppw@$      sq ~��~�c�q ~ q ~�t 983ppw@$      sq ~��~�g�q ~ q ~�t 984ppw@$      sq ~��~�kGq ~ q ~�t 985ppw@$      sq ~��~�oq ~ q ~�t 986ppw@$      sq ~��~�r�q ~ q ~�t 987ppw@$      sq ~��~�v�q ~ q ~�t 988ppw@$      sq ~��~�zKq ~ q ~�t 989ppw@$      sq ~��{b��q ~ q ~�t 99ppw@0 �s.:~sq ~��~���q ~ q ~�t 990ppw@$      sq ~��~�Тq ~ q ~�t 991ppw@$      sq ~��~��cq ~ q ~�t 992ppw@$      sq ~��~��$q ~ q ~�t 993ppw@$      sq ~��~���q ~ q ~�t 994ppw@$      sq ~��~�ߦq ~ q ~�t 995ppw@$      sq ~��~��gq ~ q ~�t 996ppw@$      sq ~��~��(q ~ q ~�t 997ppw@$      sq ~��~���q ~ q ~�t 998ppw@$      sq ~��~��q ~ q ~�t 999ppw@$      q ~��w?�      sq ~���+f3t LOGEXPt CPAPq ~��q ~ �t 0w��9�{H�sq ~���+f4q ~��q ~��q ~��q ~ �t 1w�ּ�+�y�sq ~����q ~��q ~��q ~��q ~�t 0w?�,�sq ~��K��q ~��t CPP1q ~��q ~Q�q ~=w?�IFMx[sq ~��A���q ~��q ~��q ~��q ~ �q ~Sw��,{��Wssq ~�ΐ�q ~��q ~��q ~��q ~ �q ~=w?��~0asq ~�Α���q ~��q ~��q ~��q ~ �q ~Q�w?�vN�۳sq ~�νE�,q ~��q ~��q ~��q ~ �q ~.�w?��O�b9Vsq ~������q ~��q ~��q ~��q ~ �q ~ �w��9�{H�sq ~��^~Pq ~��q ~��q ~��q ~�q ~Q�w@-��V��sq ~�ά�Lq ~��q ~��q ~��q ~�q ~ �w@Msp&��sq ~��R�NYq ~��q ~��q ~��q ~�q ~ �w@Z�LUG*sq ~��X�Irq ~��q ~��q ~��q ~WXq ~=w� �x��sq ~��ZF�5q ~��q ~��q ~��q ~WXq ~Q�w@U���"sq ~�Ψ��5q ~��q ~��q ~��q ~WXq ~ �w?�,9{t�^sq ~��d�H�q ~��q ~��q ~��q ~WXq ~�w?���>	�+sq ~�΁���q ~��q ~��q ~��q ~�q ~Sw��C���sq ~���f�Gq ~��q ~��q ~��q ~�q ~=w���ڬ��sq ~���
q ~��q ~��q ~��q ~�q ~Q�w�Ն���\�sq ~������q ~��q ~��q ~��q ~�q ~.�w��D(��W�sq ~�� c
q ~��q ~��q ~��q ~�q ~ �w����{��sq ~��ܫ��q ~��q ~��q ~��q ~�q ~�w��c3hsq ~��4Ñq ~��q ~��q ~��q ~�q ~�w?�,�sq ~��gSy"q ~��q ~��q ~��q ~�q ~ �w@�Ȭc6(sq ~��a%"�q ~��q ~��q ~��q ~�q ~�w���غ#�sq ~��1#Gq ~��q ~��q ~��q ~=q ~ �w@���u�sq ~���k�q ~��q ~��q ~��q ~=q ~�w?��=��sq ~�Ϋ8j{q ~��q ~��q ~��q ~=q ~WXw?���Y��sq ~��*��q ~��q ~��q ~��q ~=q ~�w��2�>�Asq ~��_��q ~��q ~��q ~��q ~�q ~Sw@(Ʋz2Tsq ~���j-Tq ~��q ~��q ~��q ~�q ~$�w@ �4`H�sq ~���C��q ~��q ~��q ~��q ~�q ~ �w��AL�xLsq ~��xX��q ~��q ~��q ~��q ~�q ~WXw��*�)4G�sq ~���Nbq ~��q ~��q ~��q ~�q ~�w@Y w�[sq ~��^UK�q ~��q ~��q ~��q ~�q ~hmw?�b����sq ~��d�:�q ~��q ~��q ~��q ~I�q ~WXw?���.>O�sq ~��'$�kq ~��t REPTq ~��q ~=pw�Eد�hGsq ~�����2q ~��q ~�q ~��q ~�pw��i2+csq ~��d!+�t RULEt <applypppw@�`H�sq ~����c�q ~�t <comp1pppw?�E�+�
sq ~�Ό�	�q ~�t >applypppw@FG�_��sq ~��"A�q ~�t >comp1pppw�j�^Jsq ~���کq ~�t >plural_existspppw��}���xsq ~��4::�q ~�t 	>thatlesspppw?��c�Ɩ�sq ~��Z�q ~�t >trcomp1pppw��b|�&sq ~��Կq ~�t lexpppw@J��sq ~��R롞q ~�t shift_pppppw@���λXx