�� sr -edu.cornell.cs.nlp.spf.parser.ccg.model.Model�5B��B�~ L featureSetst Ljava/util/List;L independentLexicalFeatureSetsq ~ L invalidFeaturest Ljava/util/Set;L lexicont -Ledu/cornell/cs/nlp/spf/ccg/lexicon/ILexicon;L thetat 4Ledu/cornell/cs/nlp/spf/base/hashvector/IHashVector;xpsr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.LinkedList)S]J`�"  xpw   sr Pedu.cornell.cs.nlp.spf.parser.ccg.factoredlex.features.FactoredLexicalFeatureSet�g�պ��� D 
entryScaleI lexemeNextIdD lexemeScaleI nonFactoredNextIdI templateNextIdD templateScaleL entryInitialScorert :Ledu/cornell/cs/nlp/utils/collections/ISerializableScorer;L 	lexemeIdst 5Lit/unimi/dsi/fastutil/objects/Object2IntOpenHashMap;L lexemeInitialScorerq ~ L nonFactoredIdsq ~ L templateIdsq ~ L templateInitialScorerq ~ xr Iedu.cornell.cs.nlp.spf.parser.ccg.model.lexical.AbstractLexicalFeatureSetZ���n3�� Z computeSyntaxAttributeFeaturesL 
featureTagt Ljava/lang/String;L ignoreFiltert Ljava/util/function/Predicate;xp t FACLEXsr !java.lang.invoke.SerializedLambdaoaД,)6� 
I implMethodKind[ capturedArgst [Ljava/lang/Object;L capturingClasst Ljava/lang/Class;L functionalInterfaceClassq ~ L functionalInterfaceMethodNameq ~ L "functionalInterfaceMethodSignatureq ~ L 	implClassq ~ L implMethodNameq ~ L implMethodSignatureq ~ L instantiatedMethodTypeq ~ xp   ur [Ljava.lang.Object;��X�s)l  xp    vr 0edu.cornell.cs.nlp.utils.function.PredicateUtils           xpt java/util/function/Predicatet testt (Ljava/lang/Object;)Zt 0edu/cornell/cs/nlp/utils/function/PredicateUtilst lambda$alwaysTrue$bcad8f2c$1q ~ q ~ ?�         ,?�             ?�������sr Eedu.cornell.cs.nlp.spf.parser.ccg.features.basic.scorer.UniformScorerQ�B���S D scorexp        sr 3it.unimi.dsi.fastutil.objects.Object2IntOpenHashMap         F fI sizexr 3it.unimi.dsi.fastutil.objects.AbstractObject2IntMap�o��K<z  xr 8it.unimi.dsi.fastutil.objects.AbstractObject2IntFunction�o��K<z I defRetValuexp    ?@     ,sr 9edu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.Lexeme	I����� I hashCodeCacheL 
attributesq ~ L 	constantsq ~ L 
propertiest Ljava/util/Map;L 	signaturet GLedu/cornell/cs/nlp/spf/ccg/lexicon/factored/lambda/FactoringSignature;L tokenst ,Ledu/cornell/cs/nlp/spf/base/token/TokenSeq;xp����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sr 0edu.cornell.cs.nlp.spf.mr.lambda.LogicalConstant=Q��� L baseNameq ~ L nameq ~ xr %edu.cornell.cs.nlp.spf.mr.lambda.Term�(G^� L typet .Ledu/cornell/cs/nlp/spf/mr/language/type/Type;xr 2edu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression
n�tL�h  xpsr 0edu.cornell.cs.nlp.spf.mr.language.type.TermType��6��ǭ L parentt 2Ledu/cornell/cs/nlp/spf/mr/language/type/TermType;xr ,edu.cornell.cs.nlp.spf.mr.language.type.Typeg���� I hashCodeCacheL nameq ~ xp   ct csq ~ 5  �t losq ~ 5   et ept kanpurt kanpur:cxq ~ /q ~ .sr %java.util.Collections$UnmodifiableMap��t�B L mq ~ (xpsq ~ @sr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t origint fixed_domainxsr Eedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoringSignature�ڝ�U鞉 I hashCodeI numAttributesL typesq ~ xp  E    sq ~ sr java.util.ArrayListx����a� I sizexp   w   q ~ <xq ~ Ksr *edu.cornell.cs.nlp.spf.base.token.TokenSeq�py��An I hashCode[ tokenst [Ljava/lang/String;xp�!&sur [Ljava.lang.String;��V��{G  xp   q ~ >w   
sq ~ 'A�;�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sr 3edu.cornell.cs.nlp.spf.mr.language.type.ComplexType� �g��V L domainq ~ 2L rangeq ~ 2xq ~ 7��}�t <s_pkey,<b_pkey,t>>sq ~ 5ɬ�;t s_pkeysq ~ 5 4��t pkeyq ~ <sq ~ Wq�t 
<b_pkey,t>sq ~ 5��-�t b_pkeyq ~ \sq ~ 5   tt tpt next_tot next_to:<s_pkey,<b_pkey,t>>xq ~ Uq ~ Tsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   sq ~ W?z�t 	<e,<e,t>>q ~ <sq ~ W|-t <e,t>q ~ <q ~ bxq ~ ksq ~ L��tjuq ~ O   t borderw    sq ~ '�,�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5   st sq ~ :t haryanat 	haryana:sxq ~ wq ~ vsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L)�uq ~ O   q ~ {w   sq ~ '&pxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t luckhnowt 
luckhnow:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L�<��uq ~ O   q ~ �w   +sq ~ 'QHܹsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt madhya_pradesht madhya_pradesh:sxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L�uuq ~ O   t madhyat pradeshw   sq ~ 'ȼ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt maharashtrat maharashtra:sxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L�q�uq ~ O   t theq ~ �w   !sq ~ '���ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ W��t <b_pkey,<t,s_pkey>>q ~ `sq ~ W���ot 
<t,s_pkey>q ~ bq ~ Zq ~ dt next_to:<b_pkey,<t,s_pkey>>xq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G@M�4    sq ~ sq ~ J   w   sq ~ W@M�Tt 	<e,<t,e>>q ~ <sq ~ W���t <t,e>q ~ bq ~ <xq ~ �sq ~ L���@uq ~ O   t statesw   sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t jalgaont 	jalgaon:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L���uq ~ O   q ~ �w   'sq ~ '�Ԝxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 
chandigarht chandigarh:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L|ܥuq ~ O   q ~ �w   sq ~ 'y�Ƙsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 	darbhangat darbhanga:cxq ~ �q ~ �sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~ �sq ~ L��� uq ~ O   q ~ �w   sq ~ '�I�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t kurukshetrat kurukshetra:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ LG륏uq ~ O   q ~w   $sq ~ 'R�}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t deoghart 	deoghar:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L\�2uq ~ O   q ~w   sq ~ '3>
�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt bihart bihar:sxq ~$q ~#sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~-sq ~ L�M0uq ~ O   q ~&w   sq ~ ';�Чsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~4q ~3sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~:sq ~ L;I�uq ~ O   q ~ �t statew   sq ~ 'ȆB�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~Bq ~Asq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Hsq ~ L�� puq ~ O   q ~ �w   	sq ~ '{ɡsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt 	rajasthant rajasthan:sxq ~Oq ~Nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Xsq ~ L�0��uq ~ O   q ~Qw   sq ~ '��g�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t bhusawalt 
bhusawal:cxq ~_q ~^sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~hsq ~ L䲃uq ~ O   q ~aw   sq ~ 'xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t dehradunt 
dehradun:cxq ~oq ~nsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~xsq ~ L*��uq ~ O   q ~qw   sq ~ 'PG�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t patnat patna:cxq ~q ~~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LX!�uq ~ O   q ~�w   sq ~ '�.sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�b_�uq ~ O   q ~ �q ~=t ofq ~ {w   sq ~ '�F��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t jaipurt jaipur:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�j�uq ~ O   q ~�w   )sq ~ '�^�8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t nagpurt nagpur:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�<��uq ~ O   q ~�w   sq ~ '�˴sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt 
uttrakhandt uttrakhand:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L �_tuq ~ O   q ~�w   sq ~ 'B��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt 	jharkhandt jharkhand:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lk��	uq ~ O   q ~�w   sq ~ '�|۸sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t mumbait mumbai:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L��cuq ~ O   q ~�w   #sq ~ '��h�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ yt uttar_pradesht uttar_pradesh:sxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�)�uq ~ O   t uttarq ~ �w   sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t jodhpurt 	jodhpur:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�p�"uq ~ O   q ~ w   sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t ranchit ranchi:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L��cuq ~ O   q ~w   sq ~ '�C�Xq ~Lsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ W"��nt 
<s,s_pkey>q ~ yq ~ Zt pkey_retrievert pkey_retriever:<s,s_pkey>xq ~q ~sq ~ @q ~Tsq ~ G|!<    sq ~ sq ~ J   w   sq ~ W|\t <e,e>q ~ <q ~ <xq ~&q ~Yw   sq ~ 'ڧXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t reewat reewa:cxq ~-q ~,sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~6sq ~ Lu�uq ~ O   q ~/w   sq ~ '�B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~=q ~<sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  �    sq ~ sq ~ J    w    xq ~Csq ~ L��[uq ~ O   t whichw   sq ~ '\�m�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 
aurangabadt aurangabad:cxq ~Kq ~Jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~Tsq ~ Lb+$�uq ~ O   q ~Mw   sq ~ '�Acsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t nainitalt 
nainital:cxq ~[q ~Zsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~dsq ~ Lgj(�uq ~ O   q ~]w   "sq ~ '��[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ W�!��t <b_pkey,<s_pkey,t>>q ~ `sq ~ WI�x�t 
<s_pkey,t>q ~ Zq ~ bq ~ dt next_to:<b_pkey,<s_pkey,t>>xq ~kq ~jsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ lxq ~wsq ~ L��tjuq ~ O   q ~ rw   sq ~ 'WS�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t bhopalt bhopal:cxq ~~q ~}sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�(�Puq ~ O   q ~�w   (sq ~ '�ʋq ~Lsq ~ sq ~ sq ~ 
w   q ~q ~Pxq ~�q ~�sq ~ @q ~Tsq ~ Gl�    sq ~ sq ~ J   w   q ~'q ~ <xq ~�q ~Yw   sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 	rishikesht rishikesh:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�F
uq ~ O   q ~�w   sq ~ 'H�'8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t katnit katni:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L�Wuq ~ O   q ~�w   sq ~ '\�)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Lxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ Lbau�uq ~ O   q ~ �q ~Mw   &sq ~ '��Psq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t 	mussooriet mussoorie:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L)duq ~ O   q ~�w   sq ~ 'ZR<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t gurgaont 	gurgaon:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L���uq ~ O   q ~�w   sq ~ 'Q���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t noidat noida:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ LB%�uq ~ O   q ~�w   %sq ~ '�i8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t kotat kota:cxq ~�q ~�sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~ L 2Suq ~ O   q ~�w   *sq ~ '�\�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ 8t khandwat 	khandwa:cxq ~q ~sq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~sq ~ L�=3�uq ~ O   q ~w    xsq ~ !        sq ~ #    ?@      xsq ~ #    ?@     sr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.LexicalTemplateg��%��	 I hashCodeL 	argumentsq ~ L 
propertiesq ~ (L 	signatureq ~ )L templatet 0Ledu/cornell/cs/nlp/spf/ccg/categories/Category;xp��sq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ @q ~?sq ~ G  �    sq ~ sq ~ J    w    xq ~sr 5edu.cornell.cs.nlp.spf.ccg.categories.ComplexCategory�f�Ք�nl I hashCodeCacheL syntaxt <Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/ComplexSyntax;xr .edu.cornell.cs.nlp.spf.ccg.categories.CategorycK=�.A� L 	semanticst Ljava/lang/Object;xpsr 'edu.cornell.cs.nlp.spf.mr.lambda.Lambda��Kβ�� L argumentt +Ledu/cornell/cs/nlp/spf/mr/lambda/Variable;L bodyt 4Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L typet 5Ledu/cornell/cs/nlp/spf/mr/language/type/ComplexType;xq ~ 3sr )edu.cornell.cs.nlp.spf.mr.lambda.Variable�u#$rP L 	singletonq ~ xq ~ 1q ~ <sr 5it.unimi.dsi.fastutil.objects.ReferenceSets$Singleton�7y�J| L elementq ~xpq ~'q ~'sr 4it.unimi.dsi.fastutil.objects.ReferenceSets$EmptySet�7y�J|  xpq ~'���sr :edu.cornell.cs.nlp.spf.ccg.categories.syntax.ComplexSyntax$���q\P^ I hashCodeI 	numSlahesL leftt 5Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax;L rightq ~-L slasht 4Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Slash;xr 3edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntaxʊ�	�|��  xpȠU�   sr @edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntax$SimpleSyntax��eBg� I hashCodeL 	attributeq ~ L labelq ~ xq ~/ 3�t nonet Ssq ~1 4�wq ~3t NPsr 2edu.cornell.cs.nlp.spf.ccg.categories.syntax.Slashѕ�����> C cxp /w   sq ~��sq ~ sq ~ sq ~ 
w   sq ~ 0q ~'t #0<e,e>t #0<e,e>:<e,e>xq ~<q ~;sq ~ @q ~Tsq ~ G|!<    sq ~ sq ~ J   w   q ~'xq ~Csr 4edu.cornell.cs.nlp.spf.ccg.categories.SimpleCategory��4_C� I hashCodeCacheL syntaxt BLedu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax$SimpleSyntax;xq ~sr (edu.cornell.cs.nlp.spf.mr.lambda.Literalŕtb��� [ 	argumentst 5[Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L 	predicateq ~#[ 	signaturet /[Ledu/cornell/cs/nlp/spf/mr/language/type/Type;L typeq ~ 2xq ~ 3ur 5[Ledu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression;|�㰢�[i  xp   q ~Pq ~+q ~=ur /[Ledu.cornell.cs.nlp.spf.mr.language.type.Type;>L5��  xp   q ~ <q ~ <t��Yq ~5w   sq ~��{@sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ lt #0<e,<e,t>>t #0<e,<e,t>>:<e,<e,t>>xq ~Rq ~Qsq ~ @sq ~ @sq ~ C?@     w      q ~ Eq ~ Fxsq ~ G?z��    sq ~ sq ~ J   w   q ~ lxq ~[sq ~sq ~!sq ~&q ~ <sq ~(q ~^sq ~!sq ~&q ~ <sq ~(q ~asq ~Guq ~K   q ~aq ~^sr ;it.unimi.dsi.fastutil.objects.ReferenceSets$UnmodifiableSet�7y�J|  xr Iit.unimi.dsi.fastutil.objects.ReferenceCollections$UnmodifiableCollection�7y�J| L 
collectiont 3Lit/unimi/dsi/fastutil/objects/ReferenceCollection;xpsr 2it.unimi.dsi.fastutil.objects.ReferenceOpenHashSet         F fI sizexp?@     q ~^q ~axq ~Suq ~M   q ~ <q ~ <q ~ bsq ~esq ~i?@     q ~^xq ~ nq ~+q ~ l�9��sq ~,(Iɟ   sq ~,ȠU�   q ~2q ~5sq ~7 \q ~5q ~8w   sq ~��{@sq ~ sq ~ sq ~ 
w   q ~Sxq ~tq ~ssq ~ @q ~ gsq ~ G?z��    sq ~ sq ~ J   w   q ~ lxq ~xsq ~sq ~!sq ~&q ~ <sq ~(q ~{sq ~!sq ~&q ~ <sq ~(q ~~sq ~Guq ~K   q ~{q ~~sq ~esq ~i?@     q ~~q ~{xq ~Suq ~M   q ~ <q ~ <q ~ bsq ~esq ~i?@     q ~{xq ~ nq ~+q ~ l�9��sq ~,(Iɟ   sq ~,ȠU�   q ~2q ~5q ~pq ~5q ~8w    sq ~B�V�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ <t #0et #0e:exq ~�q ~�sq ~ @q ~Tsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~Dsq ~Guq ~K   q ~�q ~+q ~uq ~M   q ~ yq ~ Z>�:q ~5w   sq ~@�H�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ @q ~Dsq ~ G  E    sq ~ sq ~ J   w   q ~ <xq ~�sq ~Dq ~�9|vq ~5w   sq ~��sq ~ sq ~ sq ~ 
w   q ~=q ~�xq ~�q ~�sq ~ @q ~Tsq ~ Gl�    sq ~ sq ~ J   w   q ~'q ~ <xq ~�sq ~Dsq ~Guq ~K   q ~�q ~+q ~=uq ~M   q ~ <q ~ <ڄs�q ~5w   sq ~��Usq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t #0<e,<t,e>>t #0<e,<t,e>>:<e,<t,e>>xq ~�q ~�sq ~ @q ~ �sq ~ G@M�4    sq ~ sq ~ J   w   q ~ �xq ~�sq ~sq ~!sq ~&q ~ nsq ~(q ~�sq ~!sq ~&q ~ <sq ~(q ~�sq ~Guq ~K   q ~�sq ~Guq ~K   q ~�sq ~esq ~i?@     q ~�q ~�xq ~�uq ~M   q ~ <q ~ bsq ~esq ~i?@     q ~�q ~�xq ~�uq ~M   q ~ <q ~ bq ~ <sq ~esq ~i?@     q ~�xq ~'q ~+sq ~ WJW'�t <<e,t>,<e,e>>q ~ nq ~'�N$!sq ~,�7�   q ~5sq ~,ȠU�   q ~2q ~5q ~pq ~8w   xsq ~ !        sr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCoordinationFeatureSet�4tHWcg+ Z cpapFeaturesZ cpp1FeaturesZ reptFeaturesxpsr Dedu.cornell.cs.nlp.spf.parser.ccg.features.basic.RuleUsageFeatureSet�k�d�L2� D scaleZ unaryRulesOnlyL 	ignoreSetq ~ xp?������� sr java.util.HashSet�D�����4  xpw   ?@      xsr Ledu.cornell.cs.nlp.spf.parser.ccg.features.basic.DynamicWordSkippingFeatures%�q�� L emptyCategoryq ~L 
featureTagq ~ xpsq ~Dp    sq ~1zT�lq ~3t EMPTYt DYNSKIPxq ~ sq ~ sq ~ J   w   q ~ xq ~�sr %java.util.Collections$UnmodifiableSet��я��U  xq ~ sq ~�w   ?@     sr .edu.cornell.cs.nlp.spf.base.hashvector.KeyArgs���]e.ɘ I hashCodeL arg1q ~ L arg2q ~ L arg3q ~ L arg4q ~ L arg5q ~ xp2Iݬq ~ t 
TMPDEFAULTpppsq ~�wzq ~ t XEMEDEFAULTpppsq ~�'��q ~ t 
LEXDEFAULTpppxsr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoredLexicon�>�"z L lexemesq ~ (L lexemesByTypeq ~ (L 	templatesq ~ (xpsq ~ C?@     0w   @   )q ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~esq ~�w   ?@     q ~Wxq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~sq ~�w   ?@     q ~xq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~{xq ~ �sq ~�w   ?@     q ~ �xq ~�sq ~�w   ?@     q ~�xq ~sq ~�w   ?@     q ~�xq ~ Nsq ~�w   ?@     q ~ +xq ~�sq ~�w   ?@     q ~�xq ~ �sq ~�w   ?@     q ~ �xq ~Isq ~�w   ?@     q ~>xq ~ �sq ~�w   ?@     q ~ �xq ~Ysq ~�w   ?@     q ~Kq ~�q ~xq ~sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~ �sq ~�w   ?@     q ~ sxq ~�sq ~�w   ?@     q ~�xq ~ �sq ~�w   ?@     q ~ �xq ~�sq ~�w   ?@     q ~�xq ~sq ~�w   ?@     q ~ xq ~.sq ~�w   ?@     q ~ xq ~Dsq ~�w   ?@     q ~9xq ~ psq ~�w   ?@     q ~ Qq ~gxq ~�sq ~�w   ?@     q ~�xq ~isq ~�w   ?@     q ~[xq ~ �sq ~�w   ?@     q ~ �xq ~7sq ~�w   ?@     q ~)xq ~ �sq ~�w   ?@     q ~ �xq ~sq ~�w   ?@     q ~
xq ~ �sq ~�w   ?@     q ~ �xq ~ysq ~�w   ?@     q ~kxq ~Usq ~�w   ?@     q ~Gxq ~;sq ~�w   ?@     q ~0xq ~�sq ~�w   ?@     q ~zxq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xxsq ~ C?@     w      q ~$sq ~�w   ?@     q ~xq ~Asq ~�w   ?@     q ~9xq ~Vsq ~�w   @?@     &q ~�q ~�q ~�q ~�q ~ �q ~�q ~zq ~�q ~0q ~
q ~Kq ~�q ~�q ~�q ~ �q ~ �q ~q ~�q ~kq ~Wq ~>q ~{q ~�q ~�q ~ q ~�q ~�q ~ �q ~ �q ~ q ~Gq ~ sq ~[q ~ �q ~ +q ~�q ~�q ~)xq ~ �sq ~�w   ?@     q ~ �xq ~�sq ~�w   ?@     q ~�xq ~ isq ~�w   ?@     q ~ Qq ~gxxsq ~ C?@     w      q ~Asq ~�w   ?@     q ~9xq ~sq ~�w   ?@     q ~xq ~�sq ~�w   ?@     q ~�q ~�xq ~�sq ~�w   ?@     q ~�xq ~�sq ~�w   ?@     q ~�xq ~vsq ~�w   ?@     q ~qq ~Oxxsr 9edu.cornell.cs.nlp.spf.base.hashvector.FastTreeHashVector;��tQ57� L valuest 0Lit/unimi/dsi/fastutil/objects/Object2DoubleMap;xpsr 5it.unimi.dsi.fastutil.objects.Object2DoubleAVLTreeMap�7y�J| I countL storedComparatort Ljava/util/Comparator;xr <it.unimi.dsi.fastutil.objects.AbstractObject2DoubleSortedMap�c����  xr 6it.unimi.dsi.fastutil.objects.AbstractObject2DoubleMap�o��K<z  xr ;it.unimi.dsi.fastutil.objects.AbstractObject2DoubleFunction�o��K<z D defRetValuexp           }psq ~�WD�t DYNSKIPppppw��      sq ~�W�"�q ~ t LEXt 0t 0pw@$      sq ~�W�"�q ~ q ~.t 0t 1pw@$      sq ~�W�&�q ~ q ~.t 1t 2pw@$      sq ~�W�i�q ~ q ~.t 10t 7pw@$      sq ~�W�m$q ~ q ~.t 11t 3pw        sq ~�W�m�q ~ q ~.t 11t 7pw@5oz�G�sq ~�W�qaq ~ q ~.t 12t 7pw@$      sq ~�W�t�q ~ q ~.t 13t 3pw        sq ~�W�u"q ~ q ~.t 13t 7pw@$      sq ~�W�xgq ~ q ~.t 14t 3pw        sq ~�W�x�q ~ q ~.t 14t 7pw@$      sq ~�W�|�q ~ q ~.t 15t 7pw@$      sq ~�W��q ~ q ~.t 16t 3pw        sq ~�WĀeq ~ q ~.t 16t 7pw@$      sq ~�Wă�q ~ q ~.t 17t 3pw        sq ~�WĄ&q ~ q ~.t 17t 7pw@F�U�i�sq ~�Wć�q ~ q ~.t 18t 7pw@$      sq ~�Wċ,q ~ q ~.t 19t 3pw        sq ~�Wċ�q ~ q ~.t 19t 7pw@$      sq ~�W�*�q ~ q ~.t 2t 3pw@$      sq ~�W�+2q ~ q ~.t 2t 7pw@$      sq ~�W��>q ~ q ~.t 20t 7pw@$      sq ~�W��q ~ q ~.t 21t 3pw        sq ~�W���q ~ q ~.t 21t 7pw@$      sq ~�W��Dq ~ q ~.t 22t 3pw        sq ~�W���q ~ q ~.t 22t 7pw@$      sq ~�W��q ~ q ~.t 23t 7pw@$      sq ~�W��Bq ~ q ~.t 24t 7pw@5oz�G�sq ~�W���q ~ q ~.t 25t 3pw        sq ~�W��q ~ q ~.t 25t 7pw@$      sq ~�W���q ~ q ~.t 26t 7pw@$      sq ~�W���q ~ q ~.t 27t 7pw@5oz�G�sq ~�W��Fq ~ q ~.t 28t 7pw@$      sq ~�W���q ~ q ~.t 29t 3pw        sq ~�W� q ~ q ~.t 29t 7pw@$      sq ~�W�.�q ~ q ~.t 3t 4pw@$      sq ~�W�R�q ~ q ~.t 30t 7pw@$      sq ~�W�U�q ~ q ~.t 31t 3pw        sq ~�W�V^q ~ q ~.t 31t 7pw@$      sq ~�W�Y�q ~ q ~.t 32t 3pw        sq ~�W�Zq ~ q ~.t 32t 7pw@$      sq ~�W�]dq ~ q ~.t 33t 3pw        sq ~�W�]�q ~ q ~.t 33t 7pw@5oz�G�sq ~�W�a%q ~ q ~.t 34t 3pw        sq ~�W�a�q ~ q ~.t 34t 7pw@$      sq ~�W�d�q ~ q ~.t 35t 3pw        sq ~�W�ebq ~ q ~.t 35t 7pw@$      sq ~�W�i#q ~ q ~.t 36t 7pw@$      sq ~�W�l�q ~ q ~.t 37t 7pw@$      sq ~�W�p)q ~ q ~.t 38t 3pw        sq ~�W�p�q ~ q ~.t 38t 7pw@5oz�G�sq ~�W�tfq ~ q ~.t 39t 7pw@$      sq ~�W�2vq ~ q ~.t 4t 5pw@$      sq ~�W�ƀq ~ q ~.t 40t 3pw        sq ~�W���q ~ q ~.t 40t 7pw@$      sq ~�W��Aq ~ q ~.t 41t 3pw        sq ~�W�ʽq ~ q ~.t 41t 7pw@$      sq ~�W��q ~ q ~.t 42t 3pw        sq ~�W��~q ~ q ~.t 42t 7pw@$      sq ~�W���q ~ q ~.t 43t 3pw        sq ~�W��?q ~ q ~.t 43t 7pw@$      sq ~�W�5�q ~ q ~.t 5t 0pw@$      sq ~�W�5�q ~ q ~.t 5t 1pw@$      sq ~�W�:q ~ q ~.t 6t 6pw@$      sq ~�W�=�q ~ q ~.t 7t 7pw@$      sq ~�W�A<q ~ q ~.t 8t 3pw        sq ~�W�A�q ~ q ~.t 8t 7pw@$      sq ~�W�D�q ~ q ~.t 9t 3pw        sq ~�W�Eyq ~ q ~.t 9t 7pw@$      q ~�w?�      sq ~�e��q ~ t TMPt 0ppw        sq ~�e���q ~ q ~�t 1ppw        sq ~�e��q ~ q ~�t 2ppw        sq ~�e�Rq ~ q ~�t 3ppw        sq ~�e�
q ~ q ~�t 4ppw        sq ~�e��q ~ q ~�t 5ppw        sq ~�e��q ~ q ~�t 6ppw        sq ~�e�Vq ~ q ~�t 7ppw        q ~�w?�      sq ~�{H�q ~ t XEMEt 0ppw@$      sq ~�{H��q ~ q ~t 1ppw@$      sq ~�{^�0q ~ q ~t 10ppw@$      sq ~�{^��q ~ q ~t 11ppw@$      sq ~�{^��q ~ q ~t 12ppw@$      sq ~�{^�sq ~ q ~t 13ppw@$      sq ~�{^�4q ~ q ~t 14ppw@$      sq ~�{_ �q ~ q ~t 15ppw@$      sq ~�{_�q ~ q ~t 16ppw@$      sq ~�{_wq ~ q ~t 17ppw@$      sq ~�{_8q ~ q ~t 18ppw@$      sq ~�{_�q ~ q ~t 19ppw@$      sq ~�{H��q ~ q ~t 2ppw@$      sq ~�{_b�q ~ q ~t 20ppw@$      sq ~�{_fPq ~ q ~t 21ppw@$      sq ~�{_jq ~ q ~t 22ppw@$      sq ~�{_m�q ~ q ~t 23ppw@$      sq ~�{_q�q ~ q ~t 24ppw@$      sq ~�{_uTq ~ q ~t 25ppw@$      sq ~�{_yq ~ q ~t 26ppw@$      sq ~�{_|�q ~ q ~t 27ppw@$      sq ~�{_��q ~ q ~t 28ppw@$      sq ~�{_�Xq ~ q ~t 29ppw@$      sq ~�{H�Dq ~ q ~t 3ppw@$      sq ~�{_��q ~ q ~t 30ppw@$      sq ~�{_گq ~ q ~t 31ppw@$      sq ~�{_�pq ~ q ~t 32ppw@$      sq ~�{_�1q ~ q ~t 33ppw@$      sq ~�{_��q ~ q ~t 34ppw@$      sq ~�{_�q ~ q ~t 35ppw@$      sq ~�{_�tq ~ q ~t 36ppw@$      sq ~�{_�5q ~ q ~t 37ppw@$      sq ~�{_��q ~ q ~t 38ppw@$      sq ~�{_��q ~ q ~t 39ppw@$      sq ~�{H�q ~ q ~t 4ppw@$      sq ~�{`KMq ~ q ~t 40ppw@$      sq ~�{`Oq ~ q ~t 41ppw@$      sq ~�{`R�q ~ q ~t 42ppw@$      sq ~�{`V�q ~ q ~t 43ppw@$      sq ~�{H��q ~ q ~t 5ppw@$      sq ~�{H��q ~ q ~t 6ppw@$      sq ~�{H�Hq ~ q ~t 7ppw@$      sq ~�{H�	q ~ q ~t 8ppw@$      sq ~�{H��q ~ q ~t 9ppw@$      q ~�w?�      x