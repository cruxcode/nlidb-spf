�� sr -edu.cornell.cs.nlp.spf.parser.ccg.model.Model�5B��B�~ L featureSetst Ljava/util/List;L independentLexicalFeatureSetsq ~ L invalidFeaturest Ljava/util/Set;L lexicont -Ledu/cornell/cs/nlp/spf/ccg/lexicon/ILexicon;L thetat 4Ledu/cornell/cs/nlp/spf/base/hashvector/IHashVector;xpsr &java.util.Collections$UnmodifiableList�%1�� L listq ~ xr ,java.util.Collections$UnmodifiableCollectionB ��^� L ct Ljava/util/Collection;xpsr java.util.LinkedList)S]J`�"  xpw   sr Pedu.cornell.cs.nlp.spf.parser.ccg.factoredlex.features.FactoredLexicalFeatureSet�g�պ��� D 
entryScaleI lexemeNextIdD lexemeScaleI nonFactoredNextIdI templateNextIdD templateScaleL entryInitialScorert :Ledu/cornell/cs/nlp/utils/collections/ISerializableScorer;L 	lexemeIdst 5Lit/unimi/dsi/fastutil/objects/Object2IntOpenHashMap;L lexemeInitialScorerq ~ L nonFactoredIdsq ~ L templateIdsq ~ L templateInitialScorerq ~ xr Iedu.cornell.cs.nlp.spf.parser.ccg.model.lexical.AbstractLexicalFeatureSetZ���n3�� Z computeSyntaxAttributeFeaturesL 
featureTagt Ljava/lang/String;L ignoreFiltert Ljava/util/function/Predicate;xp t FACLEXsr !java.lang.invoke.SerializedLambdaoaД,)6� 
I implMethodKind[ capturedArgst [Ljava/lang/Object;L capturingClasst Ljava/lang/Class;L functionalInterfaceClassq ~ L functionalInterfaceMethodNameq ~ L "functionalInterfaceMethodSignatureq ~ L 	implClassq ~ L implMethodNameq ~ L implMethodSignatureq ~ L instantiatedMethodTypeq ~ xp   ur [Ljava.lang.Object;��X�s)l  xp    vr 0edu.cornell.cs.nlp.utils.function.PredicateUtils           xpt java/util/function/Predicatet testt (Ljava/lang/Object;)Zt 0edu/cornell/cs/nlp/utils/function/PredicateUtilst lambda$alwaysTrue$bcad8f2c$1q ~ q ~ ?�        �?�             �?�������sr Eedu.cornell.cs.nlp.spf.parser.ccg.features.basic.scorer.UniformScorerQ�B���S D scorexp        sr 3it.unimi.dsi.fastutil.objects.Object2IntOpenHashMap         F fI sizexr 3it.unimi.dsi.fastutil.objects.AbstractObject2IntMap�o��K<z  xr 8it.unimi.dsi.fastutil.objects.AbstractObject2IntFunction�o��K<z I defRetValuexp    ?@    �sr 9edu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.Lexeme	I����� I hashCodeCacheL 
attributesq ~ L 	constantsq ~ L 
propertiest Ljava/util/Map;L 	signaturet GLedu/cornell/cs/nlp/spf/ccg/lexicon/factored/lambda/FactoringSignature;L tokenst ,Ledu/cornell/cs/nlp/spf/base/token/TokenSeq;xp���zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sr 0edu.cornell.cs.nlp.spf.mr.lambda.LogicalConstant=Q��� L baseNameq ~ L nameq ~ xr %edu.cornell.cs.nlp.spf.mr.lambda.Term�(G^� L typet .Ledu/cornell/cs/nlp/spf/mr/language/type/Type;xr 2edu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression
n�tL�h  xpsr 3edu.cornell.cs.nlp.spf.mr.language.type.ComplexType� �g��V L domainq ~ 2L rangeq ~ 2xr ,edu.cornell.cs.nlp.spf.mr.language.type.Typeg���� I hashCodeCacheL nameq ~ xpT��t 
<c_pkey,t>sr 0edu.cornell.cs.nlp.spf.mr.language.type.TermType��6��ǭ L parentt 2Ledu/cornell/cs/nlp/spf/mr/language/type/TermType;xq ~ 6�_Kt c_pkeysq ~ 9 4��t pkeysq ~ 9   et epsq ~ 9   tt tpt cityt city:<c_pkey,t>xq ~ /q ~ .sr %java.util.Collections$UnmodifiableMap��t�B L mq ~ (xpsq ~ Esr java.util.HashMap���`� F 
loadFactorI 	thresholdxp?@     w      t origint fixed_domainxsr Eedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoringSignature�ڝ�U鞉 I hashCodeI numAttributesL typesq ~ xp|#    sq ~ sr java.util.ArrayListx����a� I sizexp   w   sq ~ 5|-t <e,t>q ~ ?q ~ Axq ~ Psr *edu.cornell.cs.nlp.spf.base.token.TokenSeq�py��An I hashCode[ tokenst [Ljava/lang/String;xp .��ur [Ljava.lang.String;��V��{G  xp   q ~ Cw  ^sq ~ '%���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�7��t 	<i,<i,t>>sq ~ 9   it iq ~ ?sq ~ 5}�t <i,t>q ~ `q ~ At >t >:<i,<i,t>>sq ~ 0sq ~ 5I:�t 	<<e,t>,i>q ~ Qq ~ `t countt count:<<e,t>,i>sq ~ 0q ~ `t 0t 0:ixq ~ \q ~ [sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L)���    sq ~ sq ~ O   w   sq ~ 5?z�t 	<e,<e,t>>q ~ ?q ~ Qsq ~ 5I:��t 	<<e,t>,e>q ~ Qq ~ ?q ~ ?xq ~ ssq ~ S�8muq ~ V   t att leastt onew   �sq ~ 'X>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�!��t <b_pkey,<s_pkey,t>>sq ~ 9��-�t b_pkeyq ~ =sq ~ 5I�x�t 
<s_pkey,t>sq ~ 9ɬ�;t s_pkeyq ~ =q ~ At statet state:<b_pkey,<s_pkey,t>>xq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~ �sq ~ S�a�uq ~ V   t theq ~ �t ofw   �sq ~ '�˴sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 9   st ssq ~ 9  �t loq ~ ?t 
uttrakhandt uttrakhand:sxq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~ �sq ~ S �_tuq ~ V   q ~ �w  ,sq ~ 'cٔ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5l��t <lo,i>q ~ �q ~ `t sizet size:<lo,i>xq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   sq ~ 5|\t <e,e>q ~ ?q ~ ?xq ~ �sq ~ S��]uq ~ V   t smallestw   xsq ~ 'n���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5"��nt 
<s,s_pkey>q ~ �q ~ �t pkey_retrievert pkey_retriever:<s,s_pkey>xq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ �sq ~ S�� puq ~ V   t maharashtraw   �sq ~ '�݋q ~ �sq ~ sq ~ sq ~ 
w   q ~ �q ~ �xq ~ �q ~ �sq ~ Eq ~ �sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~ �q ~ �w  ysq ~ '1�̫sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5���Nt 
<c,c_pkey>sq ~ 9   ct cq ~ �q ~ ;q ~ �t pkey_retriever:<c,c_pkey>sq ~ 0q ~ �t katnit katni:cxq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~ �sq ~ S�Wuq ~ V   q ~ �w  |sq ~ '��s�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~ �sq ~ Sn�uq ~ V   t next_tow   �sq ~ ';Wvsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t haryanat 	haryana:sxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~sq ~ S�b_�uq ~ V   q ~ �q ~ �q ~ �q ~w  8sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t kanpurt kanpur:cxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~sq ~ S�!&suq ~ V   q ~w  vsq ~ 'a���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~#q ~"sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~)sq ~ S䲃uq ~ V   t bhusawalw   �sq ~ 'd�sr java.util.Collections$EmptyListz��<���  xpsq ~ sq ~ sq ~ O   w   sq ~ 0sq ~ 5T�:t 
<c_pkey,i>q ~ ;q ~ `t areat area:<c_pkey,i>xq ~2q ~1sq ~ Esq ~ Esq ~ H?@     w      q ~ Jt genlexxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~>sq ~ S�yuq ~ V   t largew  �sq ~ '�C�isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�@�t <r_pkey,<s_pkey,t>>sq ~ 9����t r_pkeyq ~ =q ~ �q ~ �t state:<r_pkey,<s_pkey,t>>xq ~Fq ~Esq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Rsq ~ S���@uq ~ V   t statesw   sq ~ 'f�g[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5\�)�t <r_pkey,<r,t>>q ~Jsq ~ 5� t <r,t>sq ~ 9   rt rq ~ �q ~ At rivert river:<r_pkey,<r,t>>xq ~Zq ~Ysq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~isq ~ S ��uq ~ V   t runw  sq ~ 'Kv/Rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5W�8dt 
<i,s_pkey>q ~ `q ~ �q ~ �t pkey_retriever:<i,s_pkey>xq ~qq ~psq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~{sq ~ S 0��uq ~ V   t havew   �sq ~ '�3� sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t uttar_pradesht uttar_pradesh:sxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�sq ~ S�)�uq ~ V   t uttart pradeshw  �sq ~ '/o��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ SȇH%uq ~ V   t riversw  ?sq ~ 'A	sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~Ht set_retrievert !set_retriever:<r_pkey,<s_pkey,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  huq ~ V   t isw  (sq ~ '� ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ tt equalst equals:<e,<e,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  huq ~ V   q ~�w   Psq ~ '�lq ~ �sq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �q ~ �t maharashtra:sxq ~�q ~�sq ~ Eq ~ �sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~ �w  usq ~ 'wѼisq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�M�
t <c_pkey,<t,s_pkey>>q ~ ;sq ~ 5���ot 
<t,s_pkey>q ~ Aq ~ �q ~ �t state:<c_pkey,<t,s_pkey>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   sq ~ 5@M�Tt 	<e,<t,e>>q ~ ?sq ~ 5���t <t,e>q ~ Aq ~ ?xq ~�sq ~ S� uq ~ V   q ~ �q ~ �w  �sq ~ '  �Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S  uq ~ V   q ~ �w   �sq ~ '��y6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5YH
t <s_pkey,<t,c_pkey>>q ~ �sq ~ 5hnI_t 
<t,c_pkey>q ~ Aq ~ ;q ~ Ct city:<s_pkey,<t,c_pkey>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S��uq ~ V   t citiesw   �sq ~ '�Ղ�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��t <t,t>q ~ Aq ~ At nott 	not:<t,t>xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~xq ~sq ~ S 3�uq ~ V   t doq ~
w   �sq ~ '�ʋsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t 	rajasthant rajasthan:sxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~"sq ~ S�0��uq ~ V   q ~w   �sq ~ '��}�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~)q ~(sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~/sq ~ SG륏uq ~ V   t kurukshetraw   sq ~ 'u\2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~ �t next_to:<s_pkey,t>xq ~7q ~6sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|#    sq ~ sq ~ O   w   q ~ Qxq ~?sq ~ Sn�uq ~ V   q ~ �w   �sq ~ '��B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5	}�Tt 
<i,c_pkey>q ~ `q ~ ;q ~ �t pkey_retriever:<i,c_pkey>xq ~Fq ~Esq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Psq ~ S ��uq ~ V   t hasw   �sq ~ 'B��isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5z���t <c_pkey,<s_pkey,t>>q ~ ;q ~ �q ~ �t state:<c_pkey,<s_pkey,t>>xq ~Xq ~Wsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~bsq ~ S� uq ~ V   q ~ �q ~ �w   ,sq ~ 'z��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~iq ~hsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~osq ~ S��cuq ~ V   t mumbaiw   ~sq ~ '^�^q ~/sq ~ sq ~ sq ~ O   w   q ~3xq ~vq ~usq ~ Eq ~9sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~zsq ~ S -��uq ~ V   q ~6w  �sq ~ 'gn8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 0��uq ~ V   q ~~w   �sq ~ ' 3~�q ~/sq ~ q ~/q ~/sq ~ Eq ~9sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S 3�uq ~ V   t manyw  �sq ~ '�)Lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ fxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~�sq ~ S 3;�uq ~ V   t mostw  +sq ~ 'OG�q ~ Ysq ~ sq ~ sq ~ 
w   q ~ ]xq ~�q ~�sq ~ Eq ~ osq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�q ~ xw   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5b?gtt <c_pkey,<c,t>>q ~ ;sq ~ 5{6ot <c,t>q ~ �q ~ Aq ~�t set_retriever:<c_pkey,<c,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  cuq ~ V   t inw  sq ~ 'z�9jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5^��pt <<e,t>,<<e,i>,e>>q ~ Qsq ~ 5H��	t 	<<e,i>,e>sq ~ 5|�t <e,i>q ~ ?q ~ `q ~ ?t argmint argmin:<<e,t>,<<e,i>,e>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   sq ~ 5W�i�t <<e,t>,<<e,e>,e>>q ~ Qsq ~ 5HgKt 	<<e,e>,e>q ~ �q ~ ?xq ~�sq ~ S��7,uq ~ V   t fewestw   asq ~ '3>
�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t bihart bihar:sxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�sq ~ S�M0uq ~ V   q ~�w  Fsq ~ 'B��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t argmaxt argmax:<<e,t>,<<e,i>,e>>q ~ fxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~�sq ~ S i�uq ~ V   q ~ �q ~�w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t ranchit ranchi:cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~sq ~ S��cuq ~ V   q ~�w   �sq ~ '�I�8q ~&sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~2t kurukshetra:cxq ~q ~
sq ~ Eq ~+sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~q ~0w  �sq ~ 'OP�rsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5"��#t 
<i,r_pkey>q ~ `q ~Jq ~ �t pkey_retriever:<i,r_pkey>xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ sq ~ S 0��uq ~ V   q ~~w   zsq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~'q ~&sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~-sq ~ S��uq ~ V   t largestw   <sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~5q ~4sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~xq ~;sq ~ S �uq ~ V   q ~
w   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5T��t 
<c_pkey,c>q ~ ;q ~ �q ~ Ct city:<c_pkey,c>xq ~Bq ~Asq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Lsq ~ S ��uq ~ V   q ~Sw   'sq ~ '��P^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5K_5�t <s_pkey,<t,i>>q ~ �sq ~ 5��it <t,i>q ~ Aq ~ `t 
populationt population:<s_pkey,<t,i>>xq ~Sq ~Rsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~`sq ~ S�b�uq ~ V   q ~Yw  ~sq ~ ' �isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5@�>t <c_pkey,s_pkey>q ~ ;q ~ �q ~ �t state:<c_pkey,s_pkey>xq ~gq ~fsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~qsq ~ S� uq ~ V   q ~ �q ~ �w   Dsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ Ct city:<c_pkey,<c,t>>xq ~xq ~wsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S ��uq ~ V   q ~Sw  )sq ~ 'm��-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S�K�uq ~ V   q ~ �q ~bw   �sq ~ '���wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5b��zt <c_pkey,<i,t>>q ~ ;q ~ bq ~�t set_retriever:<c_pkey,<i,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S ��uq ~ V   q ~Sw   �sq ~ 'u��esq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5\AV	t <r_pkey,<i,t>>q ~Jq ~ bq ~�t set_retriever:<r_pkey,<i,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 0��uq ~ V   q ~~w  $sq ~ '�?�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~�t !set_retriever:<b_pkey,<s_pkey,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  cuq ~ V   q ~�w   �sq ~ 'Q���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t noidat noida:cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�sq ~ SB%�uq ~ V   q ~�w  Ssq ~ '��,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t madhya_pradesht madhya_pradesh:sxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�sq ~ S�uuq ~ V   t madhyaq ~�w  sq ~ '�_Yq ~/sq ~ q ~/q ~/sq ~ Eq ~9sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S��uq ~ V   q ~0w  �sq ~ '��*ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5^-֟t <b_pkey,s_pkey>q ~ �q ~ �q ~ �t next_to:<b_pkey,s_pkey>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S���@uq ~ V   q ~Uw   �sq ~ '��Omsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�W	`t 
<r_pkey,r>q ~Jq ~`q ~bt river:<r_pkey,r>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	sq ~ S�K�uq ~ V   q ~ �q ~bw   5sq ~ 'ȼ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~sq ~ S�q�uq ~ V   q ~ �q ~ �w   �sq ~ '�R��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t khandwat 	khandwa:cxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~&sq ~ S�=3�uq ~ V   q ~w  �sq ~ '�89�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5KQG�t <s_pkey,<s,t>>q ~ �sq ~ 5�|_t <s,t>q ~ �q ~ Aq ~�t set_retriever:<s_pkey,<s,t>>xq ~-q ~,sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~9sq ~ S  cuq ~ V   q ~�w   �sq ~ '�C�Xq ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~?q ~>sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Cq ~#w   ]sq ~ '��q ~$sq ~ sq ~ sq ~ 
w   q ~�q ~ �xq ~Gq ~Fsq ~ Eq ~)sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~Kq ~.w  Ysq ~ '�^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5c.ͺt <c_pkey,<t,i>>q ~ ;q ~Wq ~Yt population:<c_pkey,<t,i>>xq ~Pq ~Osq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~Zsq ~ S�b�uq ~ V   q ~Yw  �sq ~ '� ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~aq ~`sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~gsq ~ S���uq ~ V   q ~ �w   �sq ~ 'E�Ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t 
aurangabadt aurangabad:cxq ~nq ~msq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~wsq ~ Sb+$�uq ~ V   q ~pw  �sq ~ '�y��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5\�Qt <r_pkey,<t,r>>q ~Jsq ~ 5���t <t,r>q ~ Aq ~`q ~bt river:<r_pkey,<t,r>>xq ~~q ~}sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ Sw�Juq ~ V   q ~bw  }sq ~ '�*�xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S 0��uq ~ V   q ~~w   6sq ~ '
wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��t <s_pkey,c_pkey>q ~ �q ~ ;q ~ �t pkey_retriever:<s_pkey,c_pkey>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  cuq ~ V   q ~�w   +sq ~ 'w#�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�sq ~ S;I�uq ~ V   q ~ �q ~ �w  �sq ~ '�Zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5c.�4t <c_pkey,<t,c>>q ~ ;sq ~ 5��t <t,c>q ~ Aq ~ �q ~ Ct city:<c_pkey,<t,c>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S .��uq ~ V   q ~ Cw   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~4q ~Yt population:<c_pkey,i>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S�yuq ~ V   q ~Aw   �sq ~ '��Zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S .��uq ~ V   q ~ Cw   0sq ~ '���9sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5I�wJt 
<s_pkey,i>q ~ �q ~ `q ~6t area:<s_pkey,i>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S 0��uq ~ V   q ~~w   �sq ~ '	�o�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5ڞJ�t <s_pkey,b_pkey>q ~ �q ~ �q ~ �t pkey_retriever:<s_pkey,b_pkey>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S  huq ~ V   q ~�w   ?sq ~ '��!�q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~q ~sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~q ~�w   �sq ~ '[�*fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~ �t next_to:<b_pkey,<s_pkey,t>>xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~ Sl	C3uq ~ V   t 	surroundsw  Isq ~ ',�?�q ~ Ysq ~ sq ~ sq ~ 
w   q ~ ]q ~ fxq ~$q ~#sq ~ Eq ~ osq ~ L�ǂ    sq ~ sq ~ O   w   q ~ tq ~ vxq ~(q ~ xw  �sq ~ '�3�`sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~-q ~,sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~3sq ~ S�p
uq ~ V   t higherw   ^sq ~ '��[�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~;q ~:sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Asq ~ S��tjuq ~ V   t borderw   �sq ~ 'E�d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �q ~oxq ~Iq ~Hsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~Osq ~ Sbau�uq ~ V   q ~ �q ~pw  �sq ~ '#:�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~Vq ~Usq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~\sq ~ S�׬�uq ~ V   t largerw  =sq ~ 'X��q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~cq ~bsq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~gq ~�w   Qsq ~ 'd��)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~Zq ~�t !set_retriever:<c_pkey,<s_pkey,t>>xq ~lq ~ksq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~tsq ~ S  huq ~ V   q ~�w  5sq ~ '�ۄ�q ~*sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~zq ~ysq ~ Eq ~/sq ~ Lo��    sq ~ sq ~ O   w   q ~ �q ~ �xq ~~q ~4w  �sq ~ ' 19�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S 0��uq ~ V   q ~~w   �sq ~ '�F��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t jaipurt jaipur:cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�sq ~ S�j�uq ~ V   q ~�w  qsq ~ '��tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  uq ~ V   q ~ �w  -sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~ �t state:<s_pkey,t>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|#    sq ~ sq ~ O   w   q ~ Qxq ~�sq ~ S���uq ~ V   q ~ �w   �sq ~ '�Gv�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S�p�"uq ~ V   t jodhpurw   Isq ~ ';�#Ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t deoghart 	deoghar:cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�sq ~ S\�2uq ~ V   q ~�w  Vsq ~ 'L>��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5J�\�t <s_pkey,<i,t>>q ~ �q ~ bq ~6t area:<s_pkey,<i,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S -��uq ~ V   q ~6w   Esq ~ 'CG�+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t gurgaont 	gurgaon:cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�sq ~ S���uq ~ V   q ~�w  nsq ~ '��I�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S0�q5uq ~ V   q ~ Ct namedq ~rw   sq ~ '�*�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ ]sq ~ 0q ~ �t 	elevationt elevation:<lo,i>xq ~	q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~sq ~ S6ǁ�uq ~ V   q ~6t thanw  sq ~ '�TP�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t nagpurt nagpur:cxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~#sq ~ S�<��uq ~ V   q ~w  %sq ~ '���,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~yxq ~*q ~)sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~0sq ~ S8~{uq ~ V   q ~ �q ~ Cq ~ �w  Xsq ~ '`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~\q ~�t set_retriever:<r_pkey,<r,t>>xq ~7q ~6sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~?sq ~ S  cuq ~ V   q ~�w  sq ~ 'm}*�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~/q ~ �t state:<s_pkey,<s,t>>xq ~Fq ~Esq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Nsq ~ S� uq ~ V   q ~ �q ~ �w   �sq ~ '*��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Uq ~Tsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~[sq ~ S:��0uq ~ V   t neighborw   �sq ~ 'N��Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ ]xq ~cq ~bsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~isq ~ S�׬�uq ~ V   q ~_w   �sq ~ 'A�;�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��}�t <s_pkey,<b_pkey,t>>q ~ �sq ~ 5q�t 
<b_pkey,t>q ~ �q ~ Aq ~ �t next_to:<s_pkey,<b_pkey,t>>xq ~pq ~osq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~|sq ~ S��tjuq ~ V   q ~Dw  dsq ~ '�T�Isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ �t state:<b_pkey,s_pkey>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S� uq ~ V   q ~ �q ~ �w   �sq ~ '�WXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S .��uq ~ V   q ~ Cw  �sq ~ 'ת��q ~`sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~�q ~�sq ~ Eq ~esq ~ Lo��    sq ~ sq ~ O   w   q ~ �q ~ �xq ~�q ~jw  �sq ~ '+u4)q ~ sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~w   sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S��5�uq ~ V   t lowestw   1sq ~ '���8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ Suq ~ V   t bordersw  sq ~ 'Y�{�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ Sn�uq ~ V   q ~ �w   Bsq ~ 'g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 0luq ~ V   t floww   �sq ~ 'xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t dehradunt 
dehradun:cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�sq ~ S*��uq ~ V   q ~�w  ]sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S  huq ~ V   q ~�w   esq ~ 'm`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~	sq ~ Sw�Juq ~ V   q ~bw   �sq ~ '�<2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ fxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~sq ~ S!N�uq ~ V   q ~ {w  Tsq ~ 'ڧXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t reewat reewa:cxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~&sq ~ Su�uq ~ V   q ~w  sq ~ 'ڿt�q ~�sq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �q ~�t 	jodhpur:cxq ~,q ~+sq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~2q ~�w  _sq ~ ' 0�nsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~7q ~6sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~=sq ~ S 0R/uq ~ V   t cant youw   dsq ~ '�ysq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Yt population:<c_pkey,<i,t>>xq ~Fq ~Esq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Nsq ~ S 0��uq ~ V   q ~~w  sq ~ 'WS�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t bhopalt bhopal:cxq ~Uq ~Tsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~^sq ~ S�(�Puq ~ V   q ~Ww  >sq ~ 'x�J�q ~ �sq ~ sq ~ sq ~ 
w   q ~�q ~ �xq ~dq ~csq ~ Eq ~ �sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~hq ~ �w  hsq ~ '!	�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Yt population:<s_pkey,i>xq ~mq ~lsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~usq ~ S�b�uq ~ V   q ~Yw   qsq ~ '��}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~|q ~{sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S 2�*uq ~ V   t livew   sq ~ 'HM�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ ]xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S�p
uq ~ V   q ~6w  Osq ~ '�&Fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5�WIt 
<r_pkey,i>q ~Jq ~ `t lengtht length:<r_pkey,i>q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Lo��    sq ~ sq ~ O   w   q ~ �q ~ �xq ~�sq ~ S��$guq ~ V   t longerw  �sq ~ ' /��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S /"�uq ~ V   t doesw   [sq ~ 't���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Qxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S 2�*uq ~ V   q ~�w  ;sq ~ '�Cdsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ fxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~�sq ~ SW��uq ~ V   q ~ �q ~ {w  Esq ~ ':�-+q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~�w  �sq ~ '
|sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  huq ~ V   q ~�w   sq ~ 'o3�dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t length:<r_pkey,<i,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S ��uq ~ V   q ~Sw   �sq ~ '�|۸q ~fsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~rt mumbai:cxq ~�q ~�sq ~ Eq ~ksq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~pw   �sq ~ '`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8xq ~ q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~ S  uq ~ V   q ~ �w   usq ~ '?�ϰsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S�;$uq ~ V   q ~�w   Usq ~ '4 2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ sq ~ SW��uq ~ V   t 	neighborsw   �sq ~ '��$�q ~�sq ~ sq ~ sq ~ 
w   q ~ fxq ~'q ~&sq ~ Eq ~�sq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~+q ~�w  'sq ~ '��P�q ~sq ~ sq ~ sq ~ 
w   q ~�xq ~/q ~.sq ~ Eq ~sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~3q ~w  &sq ~ '`6isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5|
p�t <r_pkey,s_pkey>q ~Jq ~ �q ~ �t state:<r_pkey,s_pkey>xq ~8q ~7sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Bsq ~ S���@uq ~ V   q ~Uw   sq ~ 'n��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Iq ~Hsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~Osq ~ S 3;�uq ~ V   q ~�w   tsq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ Ct 
city:<c,t>xq ~Vq ~Usq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|#    sq ~ sq ~ O   w   q ~ Qxq ~^sq ~ S .��uq ~ V   q ~ Cw  �sq ~ '�(nGsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~eq ~dsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~ksq ~ S�a�uq ~ V   t longestw  tsq ~ '{ɡq ~sq ~ sq ~ sq ~ 
w   q ~xq ~rq ~qsq ~ Eq ~sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~vq ~#w  �sq ~ '�+q ~ sq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �q ~,t 
bhusawal:cxq ~zq ~ysq ~ Eq ~%sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~*w  sq ~ '���Esq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 0��uq ~ V   q ~~w   �sq ~ '9u��q ~`sq ~ sq ~ sq ~ 
w   q ~ ]q ~�xq ~�q ~�sq ~ Eq ~esq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~�q ~jw   sq ~ 'k��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S��uq ~ V   q ~0w   �sq ~ '�\��q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~�w   Vsq ~ '�AXsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ Sgj(�uq ~ V   t nainitalw   �sq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S���uq ~ V   q ~ �w   sq ~ '�msq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S��uq ~ V   q ~0w   �sq ~ '���^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S -��uq ~ V   q ~6w   sq ~ '_�x^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~Yt population:<s_pkey,<i,t>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S�b�uq ~ V   q ~Yw   �sq ~ '|��qq ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~�w   Ssq ~ 'QHܹq ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~�w   �sq ~ '�C'�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~	q ~	sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Lo��    sq ~ sq ~ O   w   q ~ �q ~ �xq ~		sq ~ S�׬�uq ~ V   q ~_w  �sq ~ '���q ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~	q ~	sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	q ~w   ssq ~ '�u�q ~/sq ~ q ~/q ~/sq ~ Eq ~9sq ~ L  �    sq ~ sq ~ O    w    xq ~	sq ~ S�urIuq ~ V   t citizensw  �sq ~ 'eIsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~	!q ~	 sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	'sq ~ S�<��uq ~ V   t luckhnoww   sq ~ '�9�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ fxq ~	/q ~	.sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~	5sq ~ S�Xۇuq ~ V   t numberw  *sq ~ 'i�Euq ~sq ~ sq ~ sq ~ 
w   q ~
xq ~	<q ~	;sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	@q ~w   -sq ~ '^�K�q ~*sq ~ sq ~ sq ~ 
w   q ~ ]q ~�q ~�xq ~	Dq ~	Csq ~ Eq ~/sq ~ L���    sq ~ sq ~ O   w   q ~ tq ~ �q ~ �xq ~	Hq ~4w  osq ~ 'uqėsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	Mq ~	Lsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~	Ssq ~ S ��uq ~ V   q ~Sw   `sq ~ 'c�5Nq ~sq ~ sq ~ sq ~ 
w   q ~ ]q ~
q ~
xq ~	Yq ~	Xsq ~ Eq ~sq ~ L���    sq ~ sq ~ O   w   q ~ tq ~ �q ~ �xq ~	]q ~w  �sq ~ 'g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	bq ~	asq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~	hsq ~ S�+X�uq ~ V   t biggestw  sq ~ '�Q��q ~ Ysq ~ sq ~ sq ~ 
w   q ~ kxq ~	oq ~	nsq ~ Eq ~ osq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~	sq ~ xw  sq ~ '�Ӭxsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~	xq ~	wsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	~sq ~ S���uq ~ V   t jalgaonw   /sq ~ 'b�lsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t 	darbhangat darbhanga:cxq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~	�sq ~ S��� uq ~ V   q ~	�w  �sq ~ 'd��q ~�sq ~ sq ~ sq ~ 
w   q ~�q ~
xq ~	�q ~	�sq ~ Eq ~�sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~	�q ~�w  <sq ~ 'O!d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	�sq ~ S ��uq ~ V   q ~Sw   Asq ~ 'Asq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~	�sq ~ S  cuq ~ V   q ~�w   �sq ~ '���Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t 	rishikesht rishikesh:cxq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~	�sq ~ S�F
uq ~ V   q ~	�w   �sq ~ '�,�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~	�sq ~ S)�uq ~ V   q ~w  sq ~ 'gDsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~	�sq ~ S 5��uq ~ V   t runsw   csq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	�q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~	�sq ~ S��]uq ~ V   q ~ �w   sq ~ '�}8.q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~	�q ~	�sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~	�q ~�w  sq ~ 'ě}(q ~Ssq ~ sq ~ sq ~ 
w   q ~�xq ~	�q ~	�sq ~ Eq ~Xsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~	�q ~]w   �sq ~ 'X.�@sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~
 q ~	�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
sq ~ SX!�uq ~ V   t patnaw   gsq ~ '�Isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5��t <b_pkey,<t,s_pkey>>q ~ �q ~�q ~ �t state:<b_pkey,<t,s_pkey>>xq ~
q ~
sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~
sq ~ S� uq ~ V   q ~ �q ~ �w   sq ~ 'e��q ~	sq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �q ~	*t 
luckhnow:cxq ~
q ~
sq ~ Eq ~	#sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~
$q ~	(w  rsq ~ '�^�8q ~sq ~ sq ~ sq ~ 
w   q ~xq ~
(q ~
'sq ~ Eq ~sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~
,q ~$w  sq ~ '���q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~
0q ~
/sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
4q ~�w   \sq ~ 'hksq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5K_[Tt <s_pkey,<t,s>>q ~ �sq ~ 5��t <t,s>q ~ Aq ~ �q ~ �t state:<s_pkey,<t,s>>xq ~
9q ~
8sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~
Esq ~ S���@uq ~ V   q ~Uw  bsq ~ '��;Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~yxq ~
Lq ~
Ksq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~
Rsq ~ S 0��uq ~ V   q ~~w   �sq ~ '�>-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5)��t <s_pkey,r_pkey>q ~ �q ~Jq ~ �t pkey_retriever:<s_pkey,r_pkey>xq ~
Yq ~
Xsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
csq ~ S  cuq ~ V   q ~�w   �sq ~ '��3�q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~
iq ~
hsq ~ Eq ~ �sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
mq ~ �w   Zsq ~ 'z��Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~
rq ~
qsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
xsq ~ S��B"uq ~ V   t surroundingw   2sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~
�q ~
sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
�sq ~ S���uq ~ V   t 
cross_overw   �sq ~ '�.q ~ sq ~ sq ~ sq ~ 
w   q ~xq ~
�q ~
�sq ~ Eq ~sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~
�q ~w  �sq ~ '��n8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
�sq ~ Suq ~ V   q ~�w   sq ~ '�w[sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~
�sq ~ S ��uq ~ V   q ~lw  zsq ~ 'ؖE�q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~
�q ~
�sq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~
�q ~�w  `sq ~ 'R	+{sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
�sq ~ S 2Suq ~ V   t kotaw   wsq ~ 'Ԍӌq ~	�sq ~ sq ~ sq ~ 
w   q ~ �xq ~
�q ~
�sq ~ Eq ~	�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
�q ~	�w   )sq ~ 'zÛsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~
�sq ~ S��uq ~ V   t 
cross-overw  4sq ~ '�٫sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~
�sq ~ S ��uq ~ V   q ~Sw   �sq ~ 'b�/`q ~�sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~
�q ~
�sq ~ Eq ~�sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~
�q ~�w  sq ~ '��*Wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~
�sq ~ S 0��uq ~ V   q ~~w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~
�q ~
�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S 0��uq ~ V   q ~~w   7sq ~ '[
��q ~/sq ~ sq ~ sq ~ O   w   q ~3xq ~
q ~	sq ~ Eq ~9sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S��uq ~ V   q ~0w  �sq ~ '�6�Isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~ S� uq ~ V   q ~ �q ~ �w  
sq ~ 'A�r�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~"q ~!sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~(sq ~ Sz�p�uq ~ V   t sparsestw   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~0q ~/sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~6sq ~ S 2�*uq ~ V   q ~�w   �sq ~ '�Tl�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~=q ~<sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~Csq ~ S d��uq ~ V   q ~ �q ~ Cw   �sq ~ 'Lt�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Jq ~Isq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Psq ~ S ��uq ~ V   q ~Sw   Nsq ~ '1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~Wq ~Vsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~]sq ~ S���@uq ~ V   q ~Uw   �sq ~ '�U�isq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 58�3�t <r_pkey,<t,s_pkey>>q ~Jq ~�q ~ �t state:<r_pkey,<t,s_pkey>>xq ~dq ~csq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~nsq ~ S���@uq ~ V   q ~Uw  �sq ~ ':�l�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~uq ~tsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~{sq ~ Sd��Uuq ~ V   t 	excludingw   sq ~ '�� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ SĤtuq ~ V   t 	borderingw   hsq ~ '&pxq ~	sq ~ sq ~ sq ~ 
w   q ~
xq ~�q ~�sq ~ Eq ~	#sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~	(w  ksq ~ '�i8q ~
�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~
�t kota:cxq ~�q ~�sq ~ Eq ~
�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~
�w  1sq ~ '>]�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~
q ~ �t next_to:<b_pkey,<t,s_pkey>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ SW��uq ~ V   q ~#w  �sq ~ '
)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  uq ~ V   q ~ �w   {sq ~ 'IIsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~exq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S� uq ~ V   q ~ �q ~ �w  �sq ~ 'mF٦sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S���uq ~ V   q ~ �w   ksq ~ 'PG�q ~	�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~
	t patna:cxq ~�q ~�sq ~ Eq ~
sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~
w   �sq ~ '_��csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S:��0uq ~ V   q ~^w  Zsq ~ '�8��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ fxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~�sq ~ SW��uq ~ V   q ~ �q ~ {w   �sq ~ 'Z#q ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ q ~$w   sq ~ '�Оksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S ��uq ~ V   q ~Sw   Ksq ~ '{g��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5^��tt <<e,t>,<<e,i>,i>>q ~ Qsq ~ 5H���t 	<<e,i>,i>q ~�q ~ `t sumt sum:<<e,t>,<<e,i>,i>>xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~sq ~ S�ۂuq ~ V   t totalw   �sq ~ '��]sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~'q ~&sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~xq ~-sq ~ S  �uq ~ V   t now  9sq ~ '��l>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~5q ~4sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~;sq ~ S�a�uq ~ V   q ~ �q ~ �q ~ �w   Tsq ~ '�)LIsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~Bq ~Asq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Hsq ~ S� uq ~ V   q ~ �q ~ �w   Hsq ~ '  x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~Oq ~Nsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~Usq ~ S   �uq ~ V   t aw   �sq ~ '�<�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5I�x�t 
<s_pkey,s>q ~ �q ~ �q ~ �t state:<s_pkey,s>xq ~]q ~\sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~gsq ~ S���@uq ~ V   q ~Uw   "sq ~ 'XLÆq ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~mq ~lsq ~ Eq ~"sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~qq ~'w   �sq ~ '���q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~uq ~tsq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~yq ~w  �sq ~ '���hq ~`sq ~ sq ~ sq ~ 
w   q ~�xq ~}q ~|sq ~ Eq ~esq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~jw   �sq ~ '�7Tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S 5��uq ~ V   q ~	�w  isq ~ 'Q��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  uq ~ V   q ~ �w   �sq ~ 'POr�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S�~�Cuq ~ V   t combinedw  2sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S ��uq ~ V   q ~lw   
sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S ��uq ~ V   q ~Sw   �sq ~ '�89�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  huq ~ V   q ~�w   sq ~ '  ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S  �uq ~ V   t byw   �sq ~ '��w�q ~Rsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~Zsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~_w   sq ~ '�JY�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5\�/It <r_pkey,<t,i>>q ~Jq ~Wq ~�t length:<r_pkey,<t,i>>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S�;$uq ~ V   q ~�w  Gsq ~ '��&sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~sq ~ S�C�uq ~ V   t tellt mew   sq ~ 'I��q ~*sq ~ sq ~ sq ~ 
w   q ~ ]q ~�xq ~
q ~	sq ~ Eq ~/sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~q ~4w  Nsq ~ 'z�G+q ~sq ~ sq ~ sq ~ 
w   q ~ �q ~xq ~q ~sq ~ Eq ~sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~q ~w  sq ~ '	K�2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~!sq ~ SW��uq ~ V   q ~#w  csq ~ '@H�q ~Rsq ~ sq ~ sq ~ 
w   q ~ �q ~Vxq ~'q ~&sq ~ Eq ~Zsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~+q ~_w  	sq ~ '�Z�q ~ Ysq ~ sq ~ sq ~ 
w   q ~ fxq ~/q ~.sq ~ Eq ~ osq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~3q ~ xw   �sq ~ '�Z'Esq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~�t set_retriever:<s_pkey,<i,t>>xq ~8q ~7sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~@sq ~ S 0��uq ~ V   q ~~w   �sq ~ '��A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t 
chandigarht chandigarh:cxq ~Gq ~Fsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~Psq ~ S|ܥuq ~ V   q ~Iw  �sq ~ '=U5sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Wq ~Vsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~]sq ~ S6�0�uq ~ V   t highestw   �sq ~ 'OS;\q ~rsq ~ sq ~ sq ~ 
w   q ~xq ~dq ~csq ~ Eq ~wsq ~ L���    sq ~ sq ~ O   w   q ~xq ~hq ~|w  sq ~ ' �sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~mq ~lsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~ssq ~ S ��uq ~ V   t howw   �sq ~ '��usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~{q ~zsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ Sk��	uq ~ V   t 	jharkhandw   �sq ~ '��)sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S�%Cuq ~ V   t flowsw   �sq ~ 'H�'8q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~ �sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~ �w  /sq ~ 'wr�+q ~fsq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~ksq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~pw   �sq ~ '�Ԝxq ~Dsq ~ sq ~ sq ~ 
w   q ~Hxq ~�q ~�sq ~ Eq ~Lsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~Qw  esq ~ '�B�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S��[uq ~ V   t whichw   &sq ~ 'KG �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~rxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S ��uq ~ V   q ~Sw   sq ~ 'LA��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 0��uq ~ V   q ~~w   �sq ~ '��
q ~ksq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~ssq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~xw   �sq ~ '�sjIsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S� uq ~ V   q ~ �q ~ �w   sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S���uq ~ V   q ~ �w   �sq ~ '��nQq ~sq ~ sq ~ sq ~ 
w   q ~
q ~
xq ~�q ~�sq ~ Eq ~sq ~ Lo��    sq ~ sq ~ O   w   q ~ �q ~ �xq ~�q ~w  jsq ~ '���Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~q ~ sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S��uq ~ V   q ~
�w   #sq ~ 'Ojb�q ~	 sq ~ sq ~ sq ~ 
w   q ~ ]q ~�xq ~q ~sq ~ Eq ~	sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~q ~	
w  sq ~ '�Ӌ�q ~	�sq ~ sq ~ sq ~ 
w   q ~ �q ~	�xq ~q ~sq ~ Eq ~	�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~q ~	�w  �sq ~ '�8:tsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~.xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~$sq ~ S  uq ~ V   q ~ �w   �sq ~ '!�"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5Yb�,t 
<r,r_pkey>q ~`q ~Jq ~ �t pkey_retriever:<r,r_pkey>xq ~+q ~*sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~5sq ~ S  huq ~ V   q ~�w   �sq ~ '+�Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~<q ~;sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~Bsq ~ S� uq ~ V   q ~ �q ~ �w  �sq ~ '�H��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~Uq ~6t area:<s_pkey,<t,i>>xq ~Iq ~Hsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~Qsq ~ S -��uq ~ V   q ~6w  Psq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �sq ~ 0q ~ �t 	mussooriet mussoorie:cxq ~Xq ~Wsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~asq ~ S)duq ~ V   q ~Zw  wsq ~ 'W��q ~ �sq ~ sq ~ sq ~ 
w   q ~ �xq ~gq ~fsq ~ Eq ~ �sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~kq ~ �w   �sq ~ '��q ~	usq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~	�t 	jalgaon:cxq ~oq ~nsq ~ Eq ~	zsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~uq ~	w  asq ~ '�Acq ~�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~�t 
nainital:cxq ~yq ~xsq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~q ~�w  �sq ~ '�[5�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 2�*uq ~ V   q ~�w   �sq ~ '	�pIsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  uq ~ V   q ~ �w   sq ~ '-@��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S�;$uq ~ V   q ~�w  sq ~ 'i���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S6�0�uq ~ V   q ~`w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S��uq ~ V   q ~0w   ;sq ~ '�?��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S�ce|uq ~ V   t surroundw   �sq ~ '�&&>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S�a�uq ~ V   q ~ �q ~ �q ~ �w  msq ~ '�f�q ~	�sq ~ sq ~ sq ~ 
w   q ~ �q ~xq ~�q ~�sq ~ Eq ~	�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~	�w  lsq ~ ')܍�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ Sn�uq ~ V   q ~ �w  #sq ~ '�*>sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S 0luq ~ V   q ~�w   �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~ S  huq ~ V   q ~�w   Fsq ~ '%Nq ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~q ~sq ~ Eq ~"sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~q ~'w   sq ~ '�D�zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ fxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~sq ~ S c��uq ~ V   q ~vq ~�w   �sq ~ '!�"sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~$q ~#sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~*sq ~ S  cuq ~ V   q ~�w   !sq ~ '�/�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~1q ~0sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~7sq ~ S 5��uq ~ V   q ~	�w   �sq ~ '�hНsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~>q ~=sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Dsq ~ S��tjuq ~ V   q ~Dw   }sq ~ 'y�Ƙq ~	�sq ~ sq ~ sq ~ 
w   q ~	�xq ~Jq ~Isq ~ Eq ~	�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~Nq ~	�w  Hsq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Sq ~Rsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Ysq ~ S�yuq ~ V   q ~Aw   (sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~`q ~_sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~fsq ~ S�,Kuq ~ V   t withq ~ �w   sq ~ '�	��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
:xq ~nq ~msq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~tsq ~ S� uq ~ V   q ~ �q ~ �w  �sq ~ '@Z��q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~zq ~ysq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~~q ~�w   Msq ~ '�q�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ Sw�Juq ~ V   q ~bw   sq ~ '��٤sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S��aeuq ~ V   q ~�t metersw   �sq ~ '��:^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S�b�uq ~ V   q ~Yw  Rsq ~ '��q ~Dsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~Lsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~Qw   sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  cuq ~ V   q ~�w   psq ~ 'f�K�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ SȇH%uq ~ V   q ~�w   Ysq ~ '����q ~	usq ~ sq ~ sq ~ 
w   q ~ �q ~pxq ~�q ~�sq ~ Eq ~	zsq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~	w  �sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  huq ~ V   q ~�w   �sq ~ 'R�}�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~�w   �sq ~ 'L�Ӯsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ Sn�uq ~ V   q ~ �w   @sq ~ ';�t�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S���@uq ~ V   q ~Uw   �sq ~ 'Cr88sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~1q ~ �t state:<s,t>xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|#    sq ~ sq ~ O   w   q ~ Qxq ~sq ~ S���uq ~ V   q ~ �w  Dsq ~ 'ZR<�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~q ~�w   �sq ~ '�BCsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~!sq ~ S���uq ~ V   q ~
�w   �sq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~exq ~(q ~'sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~.sq ~ S���uq ~ V   q ~ �w  sq ~ '�1��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~5q ~4sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~;sq ~ S 0luq ~ V   q ~�w  ssq ~ '�7�q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~zxq ~Aq ~@sq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~Eq ~�w  �sq ~ '���Ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Jq ~Isq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Psq ~ S� uq ~ V   q ~ �q ~ �w   �sq ~ '�?��q ~&sq ~ sq ~ sq ~ 
w   q ~ �q ~xq ~Vq ~Usq ~ Eq ~+sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~Zq ~0w  Bsq ~ 'Ox��q ~�sq ~ sq ~ sq ~ 
w   q ~ ]xq ~^q ~]sq ~ Eq ~�sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~bq ~�w   Csq ~ '�*�wsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~gq ~fsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~msq ~ S ��uq ~ V   q ~Sw  0sq ~ 'ȆB�q ~ �sq ~ sq ~ sq ~ 
w   q ~�xq ~sq ~rsq ~ Eq ~ �sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~wq ~ �w   �sq ~ '��Zsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~yxq ~|q ~{sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S .��uq ~ V   q ~ Cw  Ksq ~ 'b�q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~�w   >sq ~ 'П�~q ~	�sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~	�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~	�w   �sq ~ '�x�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S���uq ~ V   q ~ �w   Rsq ~ '2�^sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~Yt population:<lo,i>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S�b�uq ~ V   q ~Yw   fsq ~ 'w�ksq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S���uq ~ V   q ~ �w  �sq ~ '~�)Usq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S��B"uq ~ V   q ~
{w  !sq ~ 'Ō�Cq ~�sq ~ sq ~ sq ~ 
w   q ~ ]q ~�q ~�xq ~�q ~�sq ~ Eq ~�sq ~ L���    sq ~ sq ~ O   w   q ~ tq ~ �q ~ �xq ~�q ~�w   �sq ~ 'eP�q ~	 sq ~ sq ~ sq ~ 
w   q ~ ]q ~�q ~�xq ~�q ~�sq ~ Eq ~	sq ~ L���    sq ~ sq ~ O   w   q ~ tq ~ �q ~ �xq ~�q ~	
w  �sq ~ '�?��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  uq ~ V   q ~ �w   �sq ~ '	�o�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  cuq ~ V   q ~�w   �sq ~ '��g�q ~ sq ~ sq ~ sq ~ 
w   q ~{xq ~�q ~�sq ~ Eq ~%sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~*w  �sq ~ ' 6�$sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~ sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~sq ~ S 6M�uq ~ V   t thatw   �sq ~ '��d�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~yxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~ S d��uq ~ V   q ~ �q ~ Cw  Qsq ~ '��y(q ~Tsq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~q ~sq ~ Eq ~Ysq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~q ~^w  7sq ~ '��q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~#q ~"sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~'q ~w   :sq ~ 'B��q ~xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �q ~�t jharkhand:sxq ~+q ~*sq ~ Eq ~}sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~1q ~�w   �sq ~ 'Q���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~6q ~5sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~<sq ~ S  cuq ~ V   q ~�w   isq ~ 'ڰ-sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Cq ~Bsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~Isq ~ S�K�uq ~ V   q ~ �q ~bw  �sq ~ '�?�	sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Pq ~Osq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Vsq ~ S  huq ~ V   q ~�w  "sq ~ '��V2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~]q ~\sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~csq ~ S 0��uq ~ V   q ~~w   sq ~ 'b�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~�q ~ Ct city:<s_pkey,c_pkey>xq ~jq ~isq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~rsq ~ S .��uq ~ V   q ~ Cw   %sq ~ '�8N[q ~Fsq ~ sq ~ sq ~ 
w   q ~ �xq ~xq ~wsq ~ Eq ~Ksq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~|q ~Pw   8sq ~ ' 1�Hsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S 1�	uq ~ V   q ~�t feetw   �sq ~ '���ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S���@uq ~ V   q ~Uw   �sq ~ ' 8)Csq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S 7�uq ~ V   q ~iw   �sq ~ '� �sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ Sn�uq ~ V   q ~ �w  fsq ~ 'f�?jsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S ��uq ~ V   q ~Sw  3sq ~ ',@b�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S�׬�uq ~ V   q ~_w  Asq ~ '~9kq ~xsq ~ sq ~ sq ~ 
w   q ~ �q ~,xq ~�q ~�sq ~ Eq ~}sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~�w  �sq ~ 'A�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  uq ~ V   q ~ �w   �sq ~ '��ژsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�q ~ fxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~�sq ~ S��7,uq ~ V   q ~�w  �sq ~ 't�7�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~^q ~bt river:<r,t>xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|#    sq ~ sq ~ O   w   q ~ Qxq ~�sq ~ Sw�Juq ~ V   q ~bw  Wsq ~ '�l
�q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~ q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~q ~�w   sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~	q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~sq ~ S6�0�uq ~ V   q ~`w   |sq ~ '�c+sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S ��uq ~ V   q ~Sw   3sq ~ '�@�gsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~#q ~"sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~)sq ~ S�@(uq ~ V   t pleasew   �sq ~ '�5�6q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~0q ~/sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~4q ~�w  sq ~ '<��6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0sq ~ 5:��t <s_pkey,<c_pkey,t>>q ~ �q ~ 7q ~ Ct city:<s_pkey,<c_pkey,t>>xq ~9q ~8sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Csq ~ S��uq ~ V   q ~w   �sq ~ '��'dsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Jq ~Isq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Psq ~ S ��uq ~ V   q ~Sw   �sq ~ 'V��q ~ Ysq ~ sq ~ sq ~ 
w   q ~ fq ~ kxq ~Vq ~Usq ~ Eq ~ osq ~ L���    sq ~ sq ~ O   w   q ~ vq ~ ?xq ~Zq ~ xw  �sq ~ '�^��q ~
�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~^q ~]sq ~ Eq ~
�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~bq ~
�w  :sq ~ '�>-�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
Zxq ~gq ~fsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~msq ~ S  huq ~ V   q ~�w   osq ~ '\�)q ~Fsq ~ sq ~ sq ~ 
w   q ~oxq ~sq ~rsq ~ Eq ~Ksq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~wq ~Pw  gsq ~ '�=�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~|q ~{sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S���uq ~ V   q ~ �w  sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S�%Cuq ~ V   q ~�w  @sq ~ '���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ SȇH%uq ~ V   q ~�w  xsq ~ 'nw4q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~�w  �sq ~ '�S�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S d��uq ~ V   q ~ �q ~ Cw   *sq ~ '��J�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~w  sq ~ 'Q���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  huq ~ V   q ~�w   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~9xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S���uq ~ V   q ~ �w    sq ~ '��\q ~sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~w  �sq ~ 'B��?q ~Fsq ~ sq ~ sq ~ 
w   q ~�q ~ fxq ~�q ~�sq ~ Eq ~Ksq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~�q ~Pw  �sq ~ '!�"�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~,xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S  uq ~ V   q ~ �w   Xsq ~ 'n�B�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�q ~�w   �sq ~ 'I �q ~ Ysq ~ sq ~ sq ~ 
w   q ~ ]q ~ kxq ~�q ~�sq ~ Eq ~ osq ~ L��S    sq ~ sq ~ O   w   q ~ tq ~ ?xq ~q ~ xw  Msq ~ 'Ғu�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~sq ~ S��tjuq ~ V   q ~Dw  .sq ~ 'z���q ~Usq ~ sq ~ sq ~ 
w   q ~ �xq ~q ~sq ~ Eq ~]sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~q ~bw   rsq ~ 'Χ�csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~qxq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~"sq ~ S:��0uq ~ V   q ~^w   �sq ~ '��3sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~)q ~(sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~/sq ~ S 0��uq ~ V   t highw   4sq ~ '}�2Csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~7q ~6sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~=sq ~ S���uq ~ V   q ~
�w   �sq ~ '����sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~Dq ~Csq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Jsq ~ SĤtuq ~ V   q ~�w   �sq ~ '���Xq ~�sq ~ sq ~ sq ~ 
w   q ~-xq ~Pq ~Osq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~Tq ~�w   msq ~ '�>.Isq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
Zxq ~Yq ~Xsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~_sq ~ S  uq ~ V   q ~ �w   Osq ~ '�2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~fq ~esq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~lsq ~ S�a�uq ~ V   q ~nw   �sq ~ '���,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Cxq ~sq ~rsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ysq ~ S8~{uq ~ V   q ~ �q ~ Cq ~ �w   Jsq ~ ')8sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ Suq ~ V   q ~�w  6sq ~ '��Qq ~/sq ~ sq ~ sq ~ O   w   q ~�q ~3xq ~�q ~�sq ~ Eq ~9sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~�q ~{w  �sq ~ '��ʉsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S���@uq ~ V   q ~Uw   �sq ~ 'l���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~[xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S�%Cuq ~ V   q ~�w   �sq ~ '9=�q ~	�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~
sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~
w   �sq ~ '^�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ Sn�uq ~ V   q ~ �w  Jsq ~ '�Jz�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ fxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~�sq ~ S i�uq ~ V   q ~ �q ~�w  Csq ~ 'L�j�q ~�sq ~ sq ~ sq ~ 
w   q ~�q ~�xq ~�q ~�sq ~ Eq ~�sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~�q ~�w   bsq ~ '�O2�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S���uq ~ V   q ~ �w  sq ~ 'h�t'q ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~�w   vsq ~ ' ��sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S z�uq ~ V   t arew   9sq ~ 'o.F-q ~sq ~ sq ~ sq ~ 
w   q ~ �xq ~�q ~�sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�q ~w   $sq ~ ' 8#Asq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~
sq ~ S 7�uq ~ V   t whatw   �sq ~ 'n�vq ~	�sq ~ sq ~ sq ~ 
w   q ~ �xq ~q ~sq ~ Eq ~	�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~q ~	�w   sq ~ '�WL�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~ sq ~ S�ce|uq ~ V   q ~�w  \sq ~ '@�eq ~�sq ~ sq ~ sq ~ 
w   q ~ �xq ~&q ~%sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~*q ~�w    sq ~ 'B�Qsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Yxq ~/q ~.sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~5sq ~ S���uq ~ V   q ~ �w  sq ~ '�\�Xq ~sq ~ sq ~ sq ~ 
w   q ~xq ~;q ~:sq ~ Eq ~"sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~?q ~'w  sq ~ 'd��$sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~mxq ~Dq ~Csq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Jsq ~ S  cuq ~ V   q ~�w   �sq ~ '&|csq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Qq ~Psq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Wsq ~ S:��0uq ~ V   q ~^w   �sq ~ '�ؿ}sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~nxq ~^q ~]sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~dsq ~ S 2�*uq ~ V   q ~�w   �sq ~ '�qRsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Gxq ~kq ~jsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~qsq ~ S 0��uq ~ V   q ~~w   nsq ~ '��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~ �xq ~xq ~wsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~~sq ~ S  uq ~ V   q ~ �w   �sq ~ 'ǥ\q ~sq ~ sq ~ sq ~ 
w   q ~ ]xq ~�q ~�sq ~ Eq ~sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�q ~w   �sq ~ '��V�q ~`sq ~ sq ~ sq ~ 
w   q ~ ]q ~�q ~�xq ~�q ~�sq ~ Eq ~esq ~ L���    sq ~ sq ~ O   w   q ~ tq ~ �q ~ �xq ~�q ~jw  [sq ~ '\�m�q ~ksq ~ sq ~ sq ~ 
w   q ~oxq ~�q ~�sq ~ Eq ~ssq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~xw  Usq ~ 'W�fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ Sl	C3uq ~ V   q ~ w   _sq ~ ' dx.sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~ S c��uq ~ V   q ~vq ~�w   Gsq ~ '�)�Vq ~�sq ~ sq ~ sq ~ 
w   q ~ ]q ~�xq ~�q ~�sq ~ Eq ~�sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~�q ~�w  sq ~ '�( ,sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S8~{uq ~ V   q ~ �q ~ Cq ~ �w  sq ~ 'oc2sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S 0��uq ~ V   q ~~w   	sq ~ '�/��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~^xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S� uq ~ V   q ~ �q ~ �w   �sq ~ '0e�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Txq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S 2�*uq ~ V   q ~�w  sq ~ 'd���sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~mxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S  uq ~ V   q ~ �w   Wsq ~ '�rSsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~ q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~ S� uq ~ V   q ~ �q ~ �w   jsq ~ '���q ~sq ~ sq ~ sq ~ 
w   q ~�q ~ fxq ~q ~sq ~ Eq ~sq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~q ~w  psq ~ ' 6Szsq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~sq ~ S 5�;uq ~ V   t showw   �sq ~ 'Ü��q ~sq ~ sq ~ sq ~ 
w   q ~ �q ~xq ~"q ~!sq ~ Eq ~"sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~&q ~'w   Lsq ~ '���Tq ~bsq ~ sq ~ sq ~ 
w   q ~�xq ~*q ~)sq ~ Eq ~gsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~.q ~lw   .sq ~ ' 8�sq ~ 
w    xsq ~ sq ~ sq ~ 
w    xq ~3q ~2sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~9sq ~ S ��uq ~ V   q ~ �w   ysq ~ '��,�q ~/sq ~ sq ~ sq ~ O   w   q ~�q ~3xq ~?q ~>sq ~ Eq ~9sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~Cq ~w  �sq ~ '`��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~8xq ~Hq ~Gsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Nsq ~ S  huq ~ V   q ~�w   sq ~ '��[Fsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~Uq ~Tsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~[sq ~ S 2ƺuq ~ V   t longw   �sq ~ ';�Чq ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~bq ~asq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~fq ~�w  Lsq ~ '���q ~/sq ~ sq ~ sq ~ O   w   q ~�sq ~ 0q ~4q ~ �t size:<c_pkey,i>xq ~jq ~isq ~ Eq ~9sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~psq ~ S�+X�uq ~ V   q ~	kw  �sq ~ '��h�q ~�sq ~ sq ~ sq ~ 
w   q ~�xq ~vq ~usq ~ Eq ~�sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~zq ~�w   �sq ~ '�>͜sq ~ 
w    xsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ At truet true:txq ~q ~~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  T    sq ~ sq ~ O   w   q ~ Axq ~�sq ~ S�Jpuq ~ V   q ~�t therew  �sq ~ '��n�q ~rsq ~ sq ~ sq ~ 
w   q ~q ~�xq ~�q ~�sq ~ Eq ~wsq ~ L�Uܘ    sq ~ sq ~ O   w   q ~q ~ txq ~�q ~|w   �sq ~ '�&��sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S�b�uq ~ V   q ~Yw   sq ~ '�Z�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~Yxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S���@uq ~ V   q ~Uw   lsq ~ '��Pq ~Usq ~ sq ~ sq ~ 
w   q ~Yxq ~�q ~�sq ~ Eq ~]sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�q ~bw  {sq ~ '�4�Xsq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~:xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~ S .��uq ~ V   q ~ Cw   sq ~ '��a�sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~
:xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S���uq ~ V   q ~ �w  �sq ~ '�<�kq ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~�w  �sq ~ '��6sq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~kxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~ S��uq ~ V   q ~w   �sq ~ '}��+q ~�sq ~ sq ~ sq ~ 
w   q ~ �q ~�xq ~�q ~�sq ~ Eq ~sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~�q ~w   =sq ~ '���ssq ~ 
w    xsq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~�sq ~ S���@uq ~ V   q ~Uw  sq ~ 'K�q ~/sq ~ sq ~ sq ~ O   w   q ~kxq ~�q ~�sq ~ Eq ~9sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~q ~qw  �sq ~ '�"l�q ~�sq ~ sq ~ sq ~ 
w   q ~�q ~
xq ~q ~sq ~ Eq ~�sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~	q ~�w  �xsq ~ !        sq ~ #    ?@      xsq ~ #    ?@     �sr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.LexicalTemplateg��%��	 I hashCodeL 	argumentsq ~ L 
propertiesq ~ (L 	signatureq ~ )L templatet 0Ledu/cornell/cs/nlp/spf/ccg/categories/Category;xpYY�Qsq ~ sq ~ sq ~ 
w   sq ~ 0q ~ vt #0<<e,t>,e>t #0<<e,t>,e>:<<e,t>,e>xq ~q ~sq ~ Eq ~sq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~sr 5edu.cornell.cs.nlp.spf.ccg.categories.ComplexCategory�f�Ք�nl I hashCodeCacheL syntaxt <Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/ComplexSyntax;xr .edu.cornell.cs.nlp.spf.ccg.categories.CategorycK=�.A� L 	semanticst Ljava/lang/Object;xpsr 'edu.cornell.cs.nlp.spf.mr.lambda.Lambda��Kβ�� L argumentt +Ledu/cornell/cs/nlp/spf/mr/lambda/Variable;L bodyt 4Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L typet 5Ledu/cornell/cs/nlp/spf/mr/language/type/ComplexType;xq ~ 3sr )edu.cornell.cs.nlp.spf.mr.lambda.Variable�u#$rP L 	singletonq ~ xq ~ 1q ~ Qsr 5it.unimi.dsi.fastutil.objects.ReferenceSets$Singleton�7y�J| L elementq ~xpq ~%sq ~sq ~$q ~ Qsq ~&q ~)sr (edu.cornell.cs.nlp.spf.mr.lambda.Literalŕtb��� [ 	argumentst 5[Ledu/cornell/cs/nlp/spf/mr/lambda/LogicalExpression;L freeVariablesq ~ L 	predicateq ~![ 	signaturet /[Ledu/cornell/cs/nlp/spf/mr/language/type/Type;L typeq ~ 2xq ~ 3ur 5[Ledu.cornell.cs.nlp.spf.mr.lambda.LogicalExpression;|�㰢�[i  xp   sq ~sq ~$q ~ ?sq ~&q ~2sq ~+uq ~/   sq ~+uq ~/   q ~2sr ;it.unimi.dsi.fastutil.objects.ReferenceSets$UnmodifiableSet�7y�J|  xr Iit.unimi.dsi.fastutil.objects.ReferenceCollections$UnmodifiableCollection�7y�J| L 
collectiont 3Lit/unimi/dsi/fastutil/objects/ReferenceCollection;xpsr 2it.unimi.dsi.fastutil.objects.ReferenceOpenHashSet         F fI sizexp?@     q ~%q ~2xq ~%ur /[Ledu.cornell.cs.nlp.spf.mr.language.type.Type;>L5��  xp   q ~ ?q ~ Asq ~+uq ~/   q ~2sq ~8sq ~<?@     q ~)q ~2xq ~)uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~%q ~)q ~2xsq ~ 0sr <edu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType&��M
� I minArgsZ orderSensitiveL optiont ELedu/cornell/cs/nlp/spf/mr/language/type/RecursiveComplexType$Option;xq ~ 5l�6�t <t*,t>q ~ Aq ~ A    sr Cedu.cornell.cs.nlp.spf.mr.language.type.RecursiveComplexType$Option�^g� �� Z isOrderSensitiveI 
minNumArgsxp    t andt 
and:<t*,t>uq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~)q ~%xq ~ Qq ~Qq ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~%xq ~ vsr 4it.unimi.dsi.fastutil.objects.ReferenceSets$EmptySet�7y�J|  xpsq ~ 5q~Et <<e,t>,<<e,t>,e>>q ~ Qq ~ vn�]sr :edu.cornell.cs.nlp.spf.ccg.categories.syntax.ComplexSyntax$���q\P^ I hashCodeI 	numSlahesL leftt 5Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax;L rightq ~[L slasht 4Ledu/cornell/cs/nlp/spf/ccg/categories/syntax/Slash;xr 3edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntaxʊ�	�|��  xp8���   sq ~Z�k�   sr @edu.cornell.cs.nlp.spf.ccg.categories.syntax.Syntax$SimpleSyntax��eBg� I hashCodeL 	attributeq ~ L labelq ~ xq ~] 3�t nonet Ssq ~ZȠU�   q ~asq ~` 4�wq ~bt NPsr 2edu.cornell.cs.nlp.spf.ccg.categories.syntax.Slashѕ�����> C cxp \sq ~g /sq ~` 3�kq ~bt Nq ~iw   �sq ~{r�|sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ �t #0<e,e>t #0<e,e>:<e,e>xq ~oq ~nsq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~vsr 4edu.cornell.cs.nlp.spf.ccg.categories.SimpleCategory��4_C� I hashCodeCacheL syntaxt BLedu/cornell/cs/nlp/spf/ccg/categories/syntax/Syntax$SimpleSyntax;xq ~sq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?4m�Pq ~ew    sq ~S	 {sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~sq ~ Eq ~"sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?GOq ~ew   ?sq ~�Yޣsq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~	�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~	�q ~Wq ~puq ~>   q ~ ?q ~ ?�Uwq ~ew   (sq ~�RVpsq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~ �sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~ �q ~Wq ~puq ~>   q ~ ?q ~ ?VM}Dq ~ew   .sq ~YE�sq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�q ~�xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~�q ~�xq ~ Qq ~�q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xnu
�sq ~Z8���   sq ~Z�f   q ~asq ~ZȠU�   q ~aq ~eq ~iq ~iq ~jq ~iw   ysq ~~W�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Eq ~�sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ vsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qsq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wsq ~ 5�~t <<<e,t>,e>,<<e,t>,e>>q ~ vq ~ v~W�!sq ~Z���z   sq ~Z�ƥ�   q ~eq ~jq ~hsq ~Z�ƥY   q ~eq ~jq ~iq ~iw   ksq ~�m��sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~	#sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~
q ~Wq ~puq ~>   q ~ ?q ~ ?�h��q ~ew   sq ~<��sq ~ sq ~ sq ~ 
w   q ~psq ~ 0q ~ �t #1<e,e>t #1<e,e>:<e,e>xq ~q ~sq ~ Eq ~	sq ~ Lo��    sq ~ sq ~ O   w   q ~ �q ~ �xq ~	sq ~sq ~sq ~$q ~ ?sq ~&q ~sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   sq ~+uq ~/   q ~q ~q ~puq ~>   q ~ ?q ~ ?sq ~+uq ~/   q ~q ~q ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~q ~xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~xq ~ Qq ~Wq ~ tBEsq ~Z�P�   sq ~` 4��q ~bt PPq ~eq ~iw   �sq ~~0�sq ~ sq ~ sq ~ 
w   q ~pxq ~$q ~#sq ~ Eq ~	�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~(sq ~wsq ~+uq ~/   q ~	�q ~Wq ~puq ~>   q ~ ?q ~ ?7+?�q ~ew   "sq ~,���sq ~ sq ~ sq ~ 
w    xq ~0q ~/sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~6sq ~sq ~sq ~$q ~ Qsq ~&q ~9sq ~sq ~$q ~ ?sq ~&q ~<sq ~+uq ~/   q ~<sq ~8sq ~<?@     q ~9q ~<xq ~9uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~9xq ~ Qq ~Wsq ~ 5JW`Lt <<e,t>,<e,t>>q ~ Qq ~ Q,���sq ~Z�9�   q ~q ~q ~iw   Rsq ~ ��sq ~ sq ~ sq ~ 
w   q ~pxq ~Kq ~Jsq ~ Eq ~isq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Osq ~sq ~sq ~$q ~ �sq ~&q ~Rsq ~sq ~$q ~ ?sq ~&q ~Usq ~+uq ~/   sq ~+uq ~/   q ~Usq ~8sq ~<?@     q ~Uq ~Rxq ~Ruq ~>   q ~ ?q ~ ?q ~[q ~puq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~Rxq ~ �q ~Wsq ~ 5�T��t <<e,e>,<e,e>>q ~ �q ~ ���=�sq ~Z�P�   q ~q ~eq ~iw   Ksq ~�x�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t #0<<e,t>,<<e,e>,e>>t %#0<<e,t>,<<e,e>,e>>:<<e,t>,<<e,e>,e>>xq ~gq ~fsq ~ Eq ~gsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~nsq ~sq ~sq ~$q ~ Qsq ~&q ~qsq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~vsq ~+uq ~/   q ~vsq ~8sq ~<?@     q ~qq ~vxq ~quq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~qxq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�q ~�q ~�uq ~>   q ~Jq ~ `q ~Wq ~�q ~}q ~huq ~>   q ~ Qq ~ �q ~ ?q ~Wq ~ v��Bsq ~Z�ƥY   q ~eq ~jq ~iw   Ysq ~V�$�sq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�q ~�q ~
uq ~>   q ~ �q ~ `q ~Wq ~�q ~�q ~huq ~>   q ~ Qq ~ �q ~ ?q ~Wq ~ v�j�sq ~Z�ƥY   q ~eq ~jq ~iw   @sq ~I�Ssq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Eq ~hsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ �sq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�xq ~ �sq ~8sq ~<?@     q ~�q ~�xq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�xq ~�q ~Wq ~��a�sq ~Z����   sq ~Z�ƥY   q ~eq ~jq ~iq ~jq ~iw   osq ~ 	��sq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~sq ~sq ~$q ~�sq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�q ~�xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~�q ~�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�q ~�q ~ �uq ~>   q ~ �q ~ `q ~Wq ~�q ~�q ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xsq ~8sq ~<?@      xsq ~ 5˹�)t <<e,i>,<<e,t>,<<e,t>,e>>>q ~�q ~X���Esq ~Z�]�   sq ~Z�ƥY   q ~eq ~jq ~iq ~q ~iw   fsq ~����sq ~ sq ~ sq ~ 
w   q ~pxq ~q ~sq ~ Eq ~]sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~wsq ~+uq ~/   q ~Yq ~Wq ~puq ~>   q ~ ?q ~ ?���q ~ew   'sq ~�;�sq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~!sq ~sq ~sq ~$q ~ Qsq ~&q ~$sq ~sq ~$q ~ Qsq ~&q ~'sq ~sq ~$q ~ ?sq ~&q ~*sq ~+uq ~/   sq ~+uq ~/   q ~*sq ~8sq ~<?@     q ~*q ~$xq ~$uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~*sq ~8sq ~<?@     q ~*q ~'xq ~'uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~*q ~$q ~'xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~$q ~'xq ~ Qsq ~8sq ~<?@     q ~$xq ~Eq ~Wsq ~ 5˪xt <<e,t>,<<e,t>,<e,t>>>q ~ Qq ~E�;�%sq ~Z8���   sq ~Z�f   q ~asq ~ZȠU�   q ~aq ~eq ~iq ~iq ~jq ~iw   >sq ~s�sq ~ sq ~ sq ~ 
w   q ~pxq ~Gq ~Fsq ~ Eq ~)sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Ksq ~sq ~sq ~$q ~ Qsq ~&q ~Nsq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~Ssq ~+uq ~/   q ~Ssq ~8sq ~<?@     q ~Sq ~Nxq ~Nuq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~Nxq ~ Qsq ~sq ~$q ~ ?sq ~&q ~]sq ~+uq ~/   q ~]q ~^q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~Zq ~�uq ~>   q ~ Qq ~�q ~ ?q ~Wq ~ v�n��sq ~Z�ƥY   q ~eq ~jq ~iw   *sq ~���sq ~ sq ~ sq ~ 
w    xq ~gq ~fsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~msq ~sq ~sq ~$q ~ Asq ~&q ~pq ~pq ~Wq ~���sq ~Z�|��   q ~aq ~aq ~iw   %sq ~�	�@sq ~ sq ~ sq ~ 
w   sq ~ 0q ~t #0<t,t>t #0<t,t>:<t,t>sq ~ 0q ~ tt #0<e,<e,t>>t #0<e,<e,t>>:<e,<e,t>>xq ~vq ~usq ~ Eq ~wsq ~ L�Uܘ    sq ~ sq ~ O   w   q ~q ~ txq ~�sq ~sq ~sq ~$q ~ ?sq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Aq ~�q ~wuq ~>   q ~ Aq ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t_p�sq ~Z�P�   q ~q ~eq ~iw   nsq ~����sq ~ sq ~ sq ~ 
w   q ~hq ~pxq ~�q ~�sq ~ Eq ~)sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~�sq ~sq ~q ~Nsq ~+uq ~/   q ~Rsq ~q ~]sq ~+uq ~/   q ~]q ~^q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~Zq ~huq ~>   q ~ Qq ~ �q ~ ?q ~Wq ~ vZ`O�q ~cw   |sq ~�գ�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~E�՟�sq ~ZmLߍ   sq ~ZȠU�   q ~aq ~eq ~hsq ~ZȠU�   q ~aq ~eq ~hq ~iw   hsq ~��sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~+sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?��|q ~ew   9sq ~W��sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?zǋq ~ew   0sq ~$/A$sq ~ sq ~ sq ~ 
w   q ~zxq ~�q ~�sq ~ Eq ~�sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~sq ~sq ~$q ~ �sq ~&q ~�sq ~sq ~$q ~Jsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�xq ~ Qsq ~8sq ~<?@     q ~�xsq ~ 5\�t <r_pkey,<e,t>>q ~Jq ~ Qq ~Wsq ~ 58-��t <<e,e>,<r_pkey,<e,t>>>q ~ �q ~�#w��sq ~Z�P�   q ~q ~eq ~iw    sq ~���Ssq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Eq ~�sq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~sq ~sq ~sq ~$q ~ Qsq ~&q ~sq ~sq ~$q ~ tsq ~&q ~	sq ~sq ~$q ~ Qsq ~&q ~sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   q ~sq ~8sq ~<?@     q ~q ~xq ~uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~ sq ~+uq ~/   sq ~+uq ~/   q ~ sq ~8sq ~<?@     q ~ q ~xq ~uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~ q ~sq ~8sq ~<?@     q ~ q ~	q ~xq ~	uq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~ q ~	q ~q ~xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~	q ~q ~xq ~ Qq ~1q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~q ~	xq ~ �sq ~8sq ~<?@     q ~q ~	q ~xq ~�uq ~>   q ~ Qq ~�q ~ ?sq ~8sq ~<?@     q ~q ~	xq ~ vsq ~8sq ~<?@     q ~xsq ~ 5�Ї�t <<e,<e,t>>,<<e,t>,e>>q ~ tq ~ vq ~Wsq ~ 5{�t <<e,t>,<<e,<e,t>>,<<e,t>,e>>>q ~ Qq ~=�
�_sq ~Z�<�   sq ~Z��;!   sq ~Z�ƥ�   q ~eq ~jq ~hsq ~Z(Iɟ   sq ~ZȠU�   q ~aq ~eq ~hq ~eq ~iq ~hq ~jq ~iw   `sq ~�L(�sq ~ sq ~ sq ~ 
w   q ~pxq ~Iq ~Hsq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Msq ~sq ~sq ~$q ~ ?sq ~&q ~Psq ~sq ~$q ~ ?sq ~&q ~Ssq ~+uq ~/   sq ~+uq ~/   q ~Sq ~Tq ~puq ~>   q ~ ?q ~ ?sq ~+uq ~/   q ~Pq ~Qq ~
uq ~>   q ~ �q ~ `sq ~8sq ~<?@     q ~Pq ~Sxq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~Pxq ~ Qq ~Wq ~ t�GOasq ~Z�P�   q ~q ~eq ~iw   sq ~x�sq ~ sq ~ sq ~ 
w    xq ~fq ~esq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~lsq ~sq ~sq ~$q ~ Qsq ~&q ~osq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~tsq ~+uq ~/   q ~tsq ~8sq ~<?@     q ~oq ~txq ~ouq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~oxq ~ Qq ~{sq ~ 0q ~ vq ~ �t the:<<e,t>,e>uq ~>   q ~ Qq ~ ?q ~Wq ~ vx~'sq ~Z�ƥY   q ~eq ~jq ~iw   bsq ~w%�bsq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Eq ~�sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ �sq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�xq ~ �q ~Wq ~aw%��sq ~Z�z�M   q ~jq ~jq ~iw   Jsq ~K��"sq ~ sq ~ sq ~ 
w   q ~wxq ~�q ~�sq ~ Eq ~7sq ~ L���    sq ~ sq ~ O   w   q ~xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Aq ~�q ~wuq ~>   q ~ Aq ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~E��sq ~Z�9�   q ~q ~q ~iw   {sq ~B�V�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ ?t #0et #0e:exq ~�q ~�sq ~ Eq ~}sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~ �uq ~>   q ~ �q ~ �>�:q ~ew   Esq ~�E�"sq ~ sq ~ sq ~ 
w   q ~wxq ~�q ~�sq ~ Eq ~)sq ~ L���    sq ~ sq ~ O   w   q ~xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Aq ~�q ~wuq ~>   q ~ Aq ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~E!d��sq ~ZmLߍ   sq ~ZȠU�   q ~aq ~eq ~hsq ~ZȠU�   q ~aq ~eq ~hq ~iw   Tsq ~���5sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Eq ~�sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ ?sq ~&q ~�q ~�q ~Wq ~ ���}Usq ~Z�|�   q ~aq ~aq ~hw   msq ~��n�sq ~ sq ~ sq ~ 
w   q ~zxq ~�q ~�sq ~ Eq ~psq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~sq ~sq ~$q ~ �sq ~&q ~�sq ~sq ~$q ~ ;sq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�xq ~ Qsq ~8sq ~<?@     q ~�xsq ~ 5b[�vt <c_pkey,<e,t>>q ~ ;q ~ Qq ~Wsq ~ 5�.�|t <<e,e>,<c_pkey,<e,t>>>q ~ �q ~
��nsq ~Z�P�   q ~q ~eq ~iw   Isq ~��{@sq ~ sq ~ sq ~ 
w   q ~zxq ~q ~sq ~ Eq ~Fsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~sq ~sq ~$q ~ ?sq ~&q ~sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   q ~q ~sq ~8sq ~<?@     q ~q ~xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~xq ~ Qq ~Wq ~ t�9��sq ~Z(Iɟ   sq ~ZȠU�   q ~aq ~eq ~hq ~eq ~iw   Vsq ~��{@sq ~ sq ~ sq ~ 
w   q ~zxq ~*q ~)sq ~ Eq ~,sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~.sq ~sq ~sq ~$q ~ ?sq ~&q ~1sq ~sq ~$q ~ ?sq ~&q ~4sq ~+uq ~/   q ~4q ~1sq ~8sq ~<?@     q ~1q ~4xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~1xq ~ Qq ~Wq ~ t�9��sq ~Z(Iɟ   sq ~ZȠU�   q ~aq ~eq ~hq ~eq ~iw   Usq ~���sq ~ sq ~ sq ~ 
w   q ~xq ~Bq ~Asq ~ Eq ~ osq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~Fsq ~sq ~sq ~$q ~ Qsq ~&q ~Isq ~sq ~$q ~ tsq ~&q ~Lsq ~sq ~$q ~ ?sq ~&q ~Osq ~+uq ~/   sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~Vsq ~+uq ~/   sq ~+uq ~/   q ~Vsq ~8sq ~<?@     q ~Iq ~Vxq ~Iuq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~Vq ~Osq ~8sq ~<?@     q ~Lq ~Vq ~Oxq ~Luq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Iq ~Lq ~Vq ~Oxq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~Iq ~Lq ~Oxq ~ Qq ~gq ~uq ~>   q ~ Qq ~ ?q ~ kq ~gq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixsq ~ 5���t <<e,<e,t>>,<e,t>>q ~ tq ~ Qq ~Wsq ~ 5�"(tt <<e,t>,<<e,<e,t>>,<e,t>>>q ~ Qq ~o	�i(sq ~Z�7F   sq ~Z��   sq ~ZȠU�   q ~aq ~eq ~hsq ~Z(Iɟ   sq ~ZȠU�   q ~aq ~eq ~hq ~eq ~iq ~hq ~jq ~iw   Xsq ~���sq ~ sq ~ sq ~ 
w   q ~pxq ~{q ~zsq ~ Eq ~Lsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~wsq ~+uq ~/   q ~Hq ~Wq ~puq ~>   q ~ ?q ~ ?E�֒q ~ew   sq ~4W��sq ~ sq ~ sq ~ 
w   q ~hq ~xq ~�q ~�sq ~ Eq ~�sq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~�sq ~sq ~q ~sq ~q ~	sq ~q ~sq ~+uq ~/   q ~sq ~q ~sq ~+uq ~/   q ~q ~1q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~q ~	xq ~ �sq ~8sq ~<?@     q ~q ~	q ~xq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~q ~	xq ~ vsq ~8sq ~<?@     q ~xq ~=q ~Wq ~?[�B�q ~Aw   �sq ~�уsq ~ sq ~ sq ~ 
w   q ~zq ~�xq ~�q ~�sq ~ Eq ~ osq ~ L��S    sq ~ sq ~ O   w   q ~ tq ~ ?xq ~�sq ~sq ~q ~Isq ~q ~Lsq ~q ~Osq ~+uq ~/   sq ~+uq ~/   q ~Uq ~gq ~ fuq ~>   q ~ Qq ~ `q ~�q ~gq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixq ~oq ~Wq ~q.r�q ~sw   ~sq ~���	sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~ �sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?Z���q ~ew   sq ~�d�sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?�{��q ~ew   /sq ~(�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Eq ~�sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~E(�>sq ~Z�|��   q ~aq ~aq ~iw   Nsq ~k�ƹsq ~ sq ~ sq ~ 
w   q ~hq ~pxq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~�sq ~sq ~sq ~$q ~ �sq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�q ~�xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~�q ~�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   q ~q ~q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~q ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xsq ~8sq ~<?@      xsq ~ 5�U�%t <<e,e>,<<e,t>,<<e,t>,e>>>q ~ �q ~X7!�sq ~Z�]�   sq ~Z�ƥY   q ~eq ~jq ~iq ~q ~iw   Asq ~
/Qsq ~ sq ~ sq ~ 
w   q ~zq ~xq ~ q ~sq ~ Eq ~�sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~$sq ~sq ~sq ~$q ~ ?sq ~&q ~'sq ~sq ~$q ~ ?sq ~&q ~*sq ~+uq ~/   sq ~+uq ~/   q ~*q ~+q ~�uq ~>   q ~Jq ~ `sq ~+uq ~/   q ~'q ~(q ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~'q ~*xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~'xq ~ Qq ~Wq ~ t�B�sq ~Z�P�   q ~q ~eq ~iw   sq ~����sq ~ sq ~ sq ~ 
w   q ~zxq ~=q ~<sq ~ Eq ~�sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~Asq ~sq ~q ~'sq ~q ~*sq ~+uq ~/   q ~.sq ~+uq ~/   q ~'q ~(q ~�uq ~>   q ~Jq ~ `sq ~8sq ~<?@     q ~'q ~*xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~'xq ~ Qq ~Wq ~ t�j<q ~9w   sq ~����sq ~ sq ~ sq ~ 
w   q ~wxq ~Rq ~Qsq ~ Eq ~wsq ~ L���    sq ~ sq ~ O   w   q ~xq ~Vsq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ ?q ~ Aq ~^q ~wuq ~>   q ~ Aq ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t ��~q ~�w   ssq ~�2.dsq ~ sq ~ sq ~ 
w   q ~hxq ~gq ~fsq ~ Eq ~	�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~ksq ~sq ~sq ~$q ~ �sq ~&q ~nsq ~sq ~$q ~ Qsq ~&q ~qsq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~vsq ~+uq ~/   q ~vsq ~8sq ~<?@     q ~vq ~qxq ~quq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~qxq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~nxq ~nuq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~nxq ~ �sq ~8sq ~<?@     q ~nq ~qxq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~nxq ~ vq ~Wsq ~ 5wй�t <<e,e>,<<e,t>,e>>q ~ �q ~ v!���sq ~Z����   sq ~Z�ƥY   q ~eq ~jq ~iq ~jq ~iw   sq ~�h��sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Eq ~5sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ ?sq ~&q ~�q ~�q ~Wq ~ ��h�sq ~Z��!�   q ~eq ~eq ~iw   csq ~оN'sq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Eq ~esq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~sq ~sq ~$q ~ ?sq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�q ~�uq ~>   q ~ �q ~ `sq ~+uq ~/   q ~�q ~�q ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t�6nzsq ~Z�P�   q ~q ~eq ~iw   
sq ~���sq ~ sq ~ sq ~ 
w   q ~zq ~xq ~�q ~�sq ~ Eq ~esq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~�sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t}6�q ~�w   �sq ~@�H�sq ~ sq ~ sq ~ 
w   q ~�xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~�sq ~wq ~�9|vq ~ew   �sq ~�
Y�sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?j�pq ~ew   sq ~��sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?t��Yq ~ew   5sq ~>�#sq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Eq ~�sq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ tsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   q ~sq ~8sq ~<?@     q ~q ~xq ~uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   sq ~+uq ~/   q ~sq ~8sq ~<?@     q ~q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~q ~sq ~8sq ~<?@     q ~q ~q ~�xq ~�uq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~q ~�q ~�q ~xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~q ~�q ~�xq ~ Qq ~&q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ �sq ~8sq ~<?@     q ~�q ~q ~�xq ~�uq ~>   q ~ Qq ~�q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ vsq ~8sq ~<?@     q ~�xq ~=q ~Wq ~?SBl/sq ~Z='S   sq ~Z�w��   sq ~Z�ƥ�   q ~eq ~jq ~hsq ~Z�P�   q ~q ~eq ~iq ~hq ~jq ~iw   �sq ~�ysq ~ sq ~ sq ~ 
w   q ~hxq ~9q ~8sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~=sq ~sq ~sq ~$q ~ Qsq ~&q ~@sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~Esq ~+uq ~/   q ~Esq ~8sq ~<?@     q ~@q ~Exq ~@uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~@xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~Osq ~+uq ~/   q ~Oq ~Pq ~�uq ~>   q ~ ;q ~ `q ~Wq ~�q ~Lq ~huq ~>   q ~ Qq ~ �q ~ ?q ~Wq ~ v>��sq ~Z�ƥY   q ~eq ~jq ~iw   asq ~IJ�sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ At #0tt #0t:txq ~Yq ~Xsq ~ Eq ~�sq ~ L  T    sq ~ sq ~ O   w   q ~ Axq ~`sq ~sq ~sq ~$q ~ ?sq ~&q ~cq ~Zsq ~8sq ~<?@      xq ~ Q
��ksq ~ZȠU�   q ~aq ~eq ~hw   �sq ~n�g@sq ~ sq ~ sq ~ 
w   q ~xq ~kq ~jsq ~ Eq ~	1sq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~osq ~sq ~sq ~$q ~ Qsq ~&q ~rsq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~wsq ~+uq ~/   q ~wsq ~8sq ~<?@     q ~rq ~wxq ~ruq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~rxq ~ Qq ~~q ~uq ~>   q ~ Qq ~ ?q ~Wq ~ v�#�Lsq ~Z�|�(   q ~aq ~jq ~iw   vsq ~��Ysq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~sq ~q ~�sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~sq ~+uq ~/   q ~q ~q ~ �uq ~>   q ~ �q ~ `q ~Wq ~�q ~q ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xsq ~8sq ~<?@      xq ~�#R�q ~w   tsq ~:��sq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Eq ~sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ tsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�q ~�xq ~�uq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�q ~�q ~�xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~�q ~�q ~�xq ~ Qq ~�q ~ fuq ~>   q ~ Qq ~ `sq ~8sq ~<?@     q ~�q ~�xq ~�sq ~8sq ~<?@     q ~�q ~�q ~�xq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ vsq ~8sq ~<?@     q ~�xq ~=q ~Wq ~?��sq ~Z='S   sq ~Z�w��   sq ~Z�ƥ�   q ~eq ~jq ~hsq ~Z�P�   q ~q ~eq ~iq ~hq ~jq ~iw   Zsq ~�[Bsq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~sq ~q ~�sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~�q ~�uq ~>   q ~ Qq ~�q ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xsq ~8sq ~<?@      xq ~˨�q ~
w   ,sq ~�x�sq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~sq ~q ~'sq ~q ~*sq ~+uq ~/   q ~.q ~1sq ~8sq ~<?@     q ~'q ~*xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~'xq ~ Qq ~Wq ~ t�A�!q ~9w   8sq ~p�sq ~ sq ~ sq ~ 
w   q ~pxq ~
q ~	sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?)�7�q ~ew   #sq ~����sq ~ sq ~ sq ~ 
w   q ~zxq ~q ~sq ~ Eq ~5sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~sq ~sq ~$q ~ �sq ~&q ~sq ~sq ~$q ~ �sq ~&q ~ sq ~sq ~$q ~ ?sq ~&q ~#sq ~+uq ~/   q ~ sq ~+uq ~/   q ~#sq ~8sq ~<?@     q ~#q ~xq ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~#q ~q ~ xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~q ~ xq ~ Qsq ~8sq ~<?@     q ~xsq ~ 5J���t <s_pkey,<e,t>>q ~ �q ~ Qq ~Wsq ~ 5�lt <<e,e>,<s_pkey,<e,t>>>q ~ �q ~3�)VNsq ~Z�P�   q ~q ~eq ~iw   <sq ~��'sq ~ sq ~ sq ~ 
w   sq ~ 0q ~ Qt #0<e,t>t #0<e,t>:<e,t>xq ~;q ~:sq ~ Eq ~ Gsq ~ L|#    sq ~ sq ~ O   w   q ~ Qxq ~Bsq ~wsq ~sq ~$q ~ ?sq ~&q ~Esq ~+uq ~/   q ~Eq ~Fq ~<uq ~>   q ~ ?q ~ Aq ~Wq ~ Q�Ǵq ~jw   [sq ~�[sq ~ sq ~ sq ~ 
w   q ~pxq ~Mq ~Lsq ~ Eq ~`sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Qsq ~sq ~sq ~$q ~ ?sq ~&q ~Tsq ~+uq ~/   q ~Tq ~Uq ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �jVB�sq ~Z��!�   q ~eq ~eq ~iw   sq ~�wK	sq ~ sq ~ sq ~ 
w   q ~pxq ~]q ~\sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~asq ~sq ~sq ~$q ~ ?sq ~&q ~dsq ~+uq ~/   q ~dq ~eq ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �jrq�sq ~Z�P�   q ~q ~eq ~iw   sq ~Q5�sq ~ sq ~ sq ~ 
w   q ~zxq ~mq ~lsq ~ Eq ~	sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~qsq ~sq ~q ~sq ~q ~sq ~+uq ~/   sq ~+uq ~/   q ~q ~q ~�uq ~>   q ~ ;q ~ `sq ~+uq ~/   q ~q ~q ~�uq ~>   q ~ ;q ~ `sq ~8sq ~<?@     q ~q ~xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~xq ~ Qq ~Wq ~ tP}sq ~w   =sq ~�K�sq ~ sq ~ sq ~ 
w   q ~zq ~pq ~xq ~�q ~�sq ~ Eq ~esq ~ L���    sq ~ sq ~ O   w   q ~ tq ~ �q ~ �xq ~�sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?sq ~+uq ~/   q ~�q ~�q ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t$��q ~�w   isq ~�3�sq ~ sq ~ sq ~ 
w   q ~zq ~pxq ~�q ~�sq ~ Eq ~/sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~�sq ~sq ~sq ~$q ~ ?sq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?sq ~+uq ~/   q ~�q ~�q ~�uq ~>   q ~ ;q ~ `sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t�^hsq ~Z�P�   q ~q ~eq ~iw   rsq ~��S7sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~Ksq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~oq ~Wq ~puq ~>   q ~ ?q ~ ?��zq ~ew   sq ~g:39sq ~ sq ~ sq ~ 
w   q ~zq ~pxq ~�q ~�sq ~ Eq ~�sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~�sq ~sq ~q ~'sq ~q ~*sq ~+uq ~/   sq ~+uq ~/   q ~*q ~+q ~puq ~>   q ~ ?q ~ ?q ~Gsq ~8sq ~<?@     q ~'q ~*xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~'xq ~ Qq ~Wq ~ t	�!q ~9w   sq ~�ҀQsq ~ sq ~ sq ~ 
w   q ~hxq ~�q ~�sq ~ Eq ~ �sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�q ~�q ~ �uq ~>   q ~ �q ~ `q ~Wq ~�q ~�q ~huq ~>   q ~ Qq ~ �q ~ ?q ~Wq ~ vdQ�sq ~Z�ƥY   q ~eq ~jq ~iw   Gsq ~1�j�sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~-q ~Wq ~puq ~>   q ~ ?q ~ ?����q ~ew   sq ~���sq ~ sq ~ sq ~ 
w    xq ~q ~sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~sq ~sq ~sq ~$q ~ Qsq ~&q ~sq ~sq ~$q ~ Qsq ~&q ~sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   sq ~+uq ~/   q ~sq ~8sq ~<?@     q ~q ~xq ~uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~sq ~8sq ~<?@     q ~q ~xq ~uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~q ~q ~xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~q ~xq ~ Qsq ~8sq ~<?@     q ~xq ~Eq ~Wq ~?���sq ~Z�g�   sq ~Z�z�z   q ~jq ~jq ~hq ~jq ~iw   esq ~��msq ~ sq ~ sq ~ 
w   q ~pxq ~0q ~/sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~4sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?|	�Aq ~ew   sq ~8/[�sq ~ sq ~ sq ~ 
w   q ~xq ~<q ~;sq ~ Eq ~sq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~@sq ~sq ~q ~�sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ �sq ~8sq ~<?@     q ~�q ~�q ~�xq ~�uq ~>   q ~ Qq ~�q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ vsq ~8sq ~<?@     q ~�xq ~=q ~Wq ~?M^�q ~�w   xsq ~G�sq ~ sq ~ sq ~ 
w   q ~xq ~Wq ~Vsq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~[sq ~sq ~q ~Psq ~q ~Ssq ~+uq ~/   sq ~+uq ~/   q ~Sq ~Tq ~
uq ~>   q ~ �q ~ `sq ~+uq ~/   q ~Pq ~Qq ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~Pq ~Sxq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~Pxq ~ Qq ~Wq ~ t�h*q ~bw   sq ~q�*�sq ~ sq ~ sq ~ 
w    xq ~oq ~nsq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~usq ~sq ~sq ~$q ~ Qsq ~&q ~xsq ~sq ~$q ~ ?sq ~&q ~{sq ~+uq ~/   q ~{sq ~8sq ~<?@     q ~xq ~{xq ~xuq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~xxq ~ Qq ~Wq ~Eq�'sq ~Z	f�   q ~sq ~ZȠU�   q ~aq ~eq ~hq ~iw   Wsq ~T��!sq ~ sq ~ sq ~ 
w   q ~zxq ~�q ~�sq ~ Eq ~ osq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~sq ~q ~Isq ~q ~Lsq ~q ~Osq ~+uq ~/   q ~�q ~ kq ~gq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixq ~oq ~Wq ~qS�0�q ~sw   $sq ~��)sq ~ sq ~ sq ~ 
w   q ~q ~�xq ~�q ~�sq ~ Eq ~ osq ~ L���    sq ~ sq ~ O   w   q ~ vq ~ ?xq ~�sq ~sq ~q ~Isq ~q ~Lsq ~q ~Osq ~+uq ~/   q ~Sq ~�q ~gq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixq ~oq ~Wq ~q��@q ~sw   �sq ~�+9Tsq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~sq ~q ~�sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~sq ~+uq ~/   q ~q ~q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~q ~�uq ~>   q ~ Qq ~�q ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xsq ~8sq ~<?@      xq ~�&`(q ~w   sq ~����sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?u��q ~ew   Msq ~�8�sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~>sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �f_hsq ~Zȡ>Z   q ~aq ~q ~iw   sq ~jw�sq ~ sq ~ sq ~ 
w   q ~zxq ~�q ~�sq ~ Eq ~sq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~�sq ~sq ~q ~Psq ~q ~Ssq ~+uq ~/   q ~aq ~Zsq ~8sq ~<?@     q ~Pq ~Sxq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Pxq ~ Qq ~Wq ~ t��q ~bw   	sq ~@#{�sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~"sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?���q ~ew   !sq ~�9Y�sq ~ sq ~ sq ~ 
w   q ~zxq ~ q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~sq ~sq ~sq ~$q ~ ?sq ~&q ~	sq ~sq ~$q ~�sq ~&q ~sq ~sq ~$q ~ ?sq ~&q ~sq ~+uq ~/   sq ~+uq ~/   q ~sq ~8sq ~<?@     q ~q ~xq ~uq ~>   q ~ ?q ~ `sq ~+uq ~/   q ~	sq ~8sq ~<?@     q ~	q ~xq ~uq ~>   q ~ ?q ~ `sq ~8sq ~<?@     q ~	q ~q ~xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~q ~	xq ~ Qsq ~8sq ~<?@     q ~	xsq ~ 5�f�At <<e,i>,<e,t>>q ~�q ~ Qq ~Wsq ~ 5���t <e,<<e,i>,<e,t>>>q ~ ?q ~$݁�sq ~Z�%   sq ~Z�P�   q ~q ~eq ~iq ~eq ~iw   sq ~n�|�sq ~ sq ~ sq ~ 
w   q ~pxq ~-q ~,sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~1sq ~sq ~q ~'sq ~q ~*sq ~+uq ~/   q ~�q ~Gsq ~8sq ~<?@     q ~'q ~*xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~'xq ~ Qq ~Wq ~ t'���q ~9w   sq ~���(sq ~ sq ~ sq ~ 
w   q ~pxq ~?q ~>sq ~ Eq ~
�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~Csq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?m��q ~ew   sq ~iQsq ~ sq ~ sq ~ 
w   q ~zq ~xq ~Kq ~Jsq ~ Eq ~ osq ~ L�ǂ    sq ~ sq ~ O   w   q ~ tq ~ vxq ~Osq ~sq ~q ~Isq ~q ~Lsq ~q ~Osq ~+uq ~/   q ~Sq ~ kq ~gq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixq ~oq ~Wq ~qhIqq ~sw   �sq ~)�Dsq ~ sq ~ sq ~ 
w   q ~zxq ~^q ~]sq ~ Eq ~Rsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~bsq ~sq ~sq ~$q ~ �sq ~&q ~esq ~sq ~$q ~ �sq ~&q ~hsq ~sq ~$q ~ ?sq ~&q ~ksq ~+uq ~/   q ~hsq ~+uq ~/   q ~ksq ~8sq ~<?@     q ~kq ~exq ~euq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~kq ~hq ~exq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~eq ~hxq ~ Qsq ~8sq ~<?@     q ~exsq ~ 5s؏�t <b_pkey,<e,t>>q ~ �q ~ Qq ~Wsq ~ 5Q3�t <<e,e>,<b_pkey,<e,t>>>q ~ �q ~{(]4�sq ~Z�P�   q ~q ~eq ~iw   sq ~D��sq ~ sq ~ sq ~ 
w   q ~zq ~pxq ~�q ~�sq ~ Eq ~esq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~�sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?sq ~+uq ~/   q ~�q ~�q ~�uq ~>   q ~ �q ~ `sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t�ٱ�q ~�w   }sq ~�P3�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�q ~�q ~�xq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~�q ~�xq ~ Qsq ~8sq ~<?@     q ~�xq ~Eq ~Wq ~?�P/�sq ~Z8���   sq ~Z�k�   q ~asq ~ZȠU�   q ~aq ~eq ~hq ~iq ~jq ~iw   sq ~��o�sq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~	�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?@��q ~ew   Bsq ~�7�msq ~ sq ~ sq ~ 
w   q ~pxq ~�q ~�sq ~ Eq ~
sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?;2�Aq ~ew   sq ~Ɓgsq ~ sq ~ sq ~ 
w   q ~xq ~�q ~�sq ~ Eq ~/sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~�sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�q ~�uq ~>   q ~ ;q ~ `sq ~+uq ~/   q ~�q ~�q ~uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t�>��q ~�w   4sq ~��v�sq ~ sq ~ sq ~ 
w    xq ~�q ~�sq ~ Eq ~�sq ~ L  �    sq ~ sq ~ O    w    xq ~�sq ~sq ~sq ~$q ~ Qsq ~&q ~�sq ~sq ~$q ~ ?sq ~&q ~�sq ~+uq ~/   q ~�sq ~8sq ~<?@     q ~�q ~�xq ~�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~E��r�sq ~Z(J�]   sq ~ZȠU�   q ~aq ~eq ~hq ~q ~iw   sq ~GsJ�sq ~ sq ~ sq ~ 
w   q ~wxq ~ q ~ sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L���    sq ~ sq ~ O   w   q ~xq ~ sq ~sq ~sq ~$q ~ Qsq ~&q ~ sq ~sq ~$q ~ ?sq ~&q ~ sq ~+uq ~/   sq ~+uq ~/   q ~ sq ~8sq ~<?@     q ~ q ~ xq ~ uq ~>   q ~ ?q ~ Aq ~ q ~wuq ~>   q ~ Aq ~ Asq ~8sq ~<?@     q ~ xq ~ Qq ~Wq ~E|�[�sq ~Z�z�M   q ~jq ~jq ~iw   ^sq ~ܞf�sq ~ sq ~ sq ~ 
w   q ~pxq ~ )q ~ (sq ~ Eq ~%sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ -sq ~wsq ~+uq ~/   q ~{q ~Wq ~puq ~>   q ~ ?q ~ ?���pq ~ew   sq ~f{!sq ~ sq ~ sq ~ 
w   q ~pxq ~ 5q ~ 4sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ 9sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?vG�q ~ew   2sq ~q�%{sq ~ sq ~ sq ~ 
w    xq ~ Aq ~ @sq ~ Eq ~sq ~ L  �    sq ~ sq ~ O    w    xq ~ Esq ~sq ~sq ~$q ~ Qsq ~&q ~ Hsq ~sq ~$q ~ ?sq ~&q ~ Ksq ~+uq ~/   q ~ Ksq ~8sq ~<?@     q ~ Kq ~ Hxq ~ Huq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~ Hxq ~ Qq ~Wq ~Eq�!�sq ~Z	aJ   q ~sq ~ZȠU�   q ~aq ~eq ~iq ~iw   dsq ~)U$�sq ~ sq ~ sq ~ 
w   q ~pxq ~ Yq ~ Xsq ~ Eq ~Zsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ ]sq ~wsq ~+uq ~/   q ~Vq ~Wq ~puq ~>   q ~ ?q ~ ?�PK�q ~ew   sq ~�y��sq ~ sq ~ sq ~ 
w   q ~hxq ~ eq ~ dsq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~ isq ~sq ~sq ~$q ~ �sq ~&q ~ lsq ~sq ~$q ~ Qsq ~&q ~ osq ~sq ~$q ~ Qsq ~&q ~ rsq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~ wsq ~+uq ~/   sq ~+uq ~/   q ~ wsq ~8sq ~<?@     q ~ wq ~ oxq ~ ouq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~ wsq ~8sq ~<?@     q ~ wq ~ rxq ~ ruq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~ wq ~ rq ~ oxq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~ rq ~ oxq ~ Qsq ~sq ~$q ~ ?sq ~&q ~ �sq ~+uq ~/   q ~ �sq ~8sq ~<?@     q ~ �q ~ lxq ~ luq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~ lxq ~ �sq ~8sq ~<?@     q ~ rq ~ lq ~ oxq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~ lq ~ oxq ~ vsq ~8sq ~<?@     q ~ lxq ~Xq ~Wq ~\�sq ~Z(��O   sq ~Z�]�   sq ~Z�ƥY   q ~eq ~jq ~iq ~q ~iq ~jq ~iw   Lsq ~��B�sq ~ sq ~ sq ~ 
w   q ~zq ~q ~�xq ~ �q ~ �sq ~ Eq ~ osq ~ L)���    sq ~ sq ~ O   w   q ~ tq ~ vq ~ ?xq ~ �sq ~sq ~q ~Isq ~q ~Lsq ~q ~Osq ~+uq ~/   sq ~+uq ~/   q ~Uq ~gq ~uq ~>   q ~ Qq ~ ?q ~�q ~gq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixq ~oq ~Wq ~qB��q ~sw   lsq ~���^sq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~ �sq ~sq ~sq ~$q ~ Qsq ~&q ~ �sq ~sq ~$q ~ ?sq ~&q ~ �sq ~+uq ~/   q ~ �sq ~8sq ~<?@     q ~ �q ~ �xq ~ �uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~ �xq ~ Qq ~Wq ~E���~sq ~ZmL1-   sq ~ZȠU�   q ~aq ~eq ~isq ~ZȠU�   q ~aq ~eq ~iq ~iw   3sq ~n@��sq ~ sq ~ sq ~ 
w   q ~pxq ~ �q ~ �sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ �sq ~wsq ~+uq ~/   q ~zq ~Wq ~puq ~>   q ~ ?q ~ ?';�Yq ~ew   &sq ~K�=sq ~ sq ~ sq ~ 
w   q ~pxq ~ �q ~ �sq ~ Eq ~esq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~ �sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t�?q ~�w   )sq ~(W~sq ~ sq ~ sq ~ 
w    xq ~ �q ~ �sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~ �sq ~sq ~sq ~$q ~ Qsq ~&q ~ �sq ~sq ~$q ~ ?sq ~&q ~ �sq ~+uq ~/   q ~ �sq ~8sq ~<?@     q ~ �q ~ �xq ~ �uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~ �xq ~ Qq ~Wq ~E(S�sq ~Z�z�M   q ~jq ~jq ~iw   Ssq ~��2"sq ~ sq ~ sq ~ 
w   q ~pxq ~!	q ~!sq ~ Eq ~}sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~!sq ~wsq ~+uq ~/   q ~,q ~Wq ~puq ~>   q ~ ?q ~ ?U�X�q ~ew   sq ~Ïn�sq ~ sq ~ sq ~ 
w   q ~hq ~xq ~!q ~!sq ~ Eq ~sq ~ L���    sq ~ sq ~ O   w   q ~�q ~ vxq ~!sq ~sq ~q ~�sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ �sq ~8sq ~<?@     q ~�q ~�q ~�xq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�q ~�xq ~ vsq ~8sq ~<?@     q ~�xq ~=q ~Wq ~?�.-�q ~�w   _sq ~G0�Hsq ~ sq ~ sq ~ 
w   q ~zxq ~!0q ~!/sq ~ Eq ~wsq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~!4sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Aq ~!<q ~uq ~>   q ~ Aq ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ tFx��q ~�w   :sq ~�^�sq ~ sq ~ sq ~ 
w   q ~�xq ~!Eq ~!Dsq ~ Eq ~ osq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~!Isq ~sq ~q ~Isq ~q ~Lsq ~q ~Osq ~+uq ~/   q ~�q ~�q ~gq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~Lq ~Ixq ~ Qsq ~8sq ~<?@     q ~Ixq ~oq ~Wq ~q���|q ~sw   Osq ~�H��sq ~ sq ~ sq ~ 
w   q ~pxq ~!Xq ~!Wsq ~ Eq ~	zsq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~!\sq ~wsq ~+uq ~/   q ~pq ~Wq ~puq ~>   q ~ ?q ~ ?�C�yq ~ew   Fsq ~��p�sq ~ sq ~ sq ~ 
w   q ~xq ~!dq ~!csq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ LI:�t    sq ~ sq ~ O   w   q ~ vxq ~!jsq ~sq ~sq ~$q ~ Qsq ~&q ~!msq ~sq ~$q ~ tsq ~&q ~!psq ~sq ~$q ~ Qsq ~&q ~!ssq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~!xsq ~+uq ~/   q ~!xsq ~8sq ~<?@     q ~!xq ~!sxq ~!suq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~!sxq ~ Qsq ~sq ~$q ~ ?sq ~&q ~!�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~!�sq ~+uq ~/   sq ~+uq ~/   q ~!�sq ~8sq ~<?@     q ~!�q ~!mxq ~!muq ~>   q ~ ?q ~ Asq ~+uq ~/   q ~!�q ~!�sq ~8sq ~<?@     q ~!�q ~!�q ~!pxq ~!puq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~!�q ~!�q ~!pq ~!mxq ~Guq ~>   q ~ Aq ~ Aq ~ Asq ~8sq ~<?@     q ~!pq ~!�q ~!mxq ~ Qq ~!�q ~uq ~>   q ~ Qq ~ ?sq ~8sq ~<?@     q ~!mq ~!pxq ~ �sq ~8sq ~<?@     q ~!pq ~!sq ~!mxq ~�uq ~>   q ~ Qq ~�q ~ ?sq ~8sq ~<?@     q ~!mq ~!pxq ~ vsq ~8sq ~<?@     q ~!mxq ~=q ~Wq ~?�&��sq ~Z�<�   sq ~Z��;!   sq ~Z�ƥ�   q ~eq ~jq ~hsq ~Z(Iɟ   sq ~ZȠU�   q ~aq ~eq ~hq ~eq ~iq ~hq ~jq ~iw   wsq ~	7�sq ~ sq ~ sq ~ 
w   q ~zq ~xq ~!�q ~!�sq ~ Eq ~	sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~!�sq ~sq ~q ~sq ~q ~sq ~+uq ~/   q ~wq ~sq ~8sq ~<?@     q ~q ~xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~xq ~ Qq ~Wq ~ t�?Qq ~w   usq ~rS{�sq ~ sq ~ sq ~ 
w   q ~pxq ~!�q ~!�sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~!�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?+N��q ~ew   7sq ~l�b�sq ~ sq ~ sq ~ 
w   q ~pxq ~!�q ~!�sq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~!�sq ~wsq ~+uq ~/   q ~q ~Wq ~puq ~>   q ~ ?q ~ ?%��`q ~ew   Qsq ~ʆ�sq ~ sq ~ sq ~ 
w   q ~zq ~pxq ~!�q ~!�sq ~ Eq ~sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~!�sq ~sq ~q ~Psq ~q ~Ssq ~+uq ~/   q ~Wq ~Zsq ~8sq ~<?@     q ~Pq ~Sxq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Pxq ~ Qq ~Wq ~ tmG��q ~bw   �sq ~���sq ~ sq ~ sq ~ 
w    xq ~!�q ~!�sq ~ Esq ~ Esq ~ H?@     w      q ~ Jq ~ Kxsq ~ L  �    sq ~ sq ~ O    w    xq ~!�sq ~sq ~sq ~$q ~ Asq ~&q ~!�q ~!�q ~Wq ~���sq ~Z�|�   q ~aq ~aq ~hw   jsq ~��sq ~ sq ~ sq ~ 
w    xq ~!�q ~!�sq ~ Eq ~�sq ~ L  �    sq ~ sq ~ O    w    xq ~!�sq ~sq ~sq ~$q ~ ?sq ~&q ~!�q ~!�q ~Wq ~ ����sq ~ZȠU�   q ~aq ~eq ~iw   ]sq ~(�Ysq ~ sq ~ sq ~ 
w    xq ~"q ~"sq ~ Eq ~sq ~ L  �    sq ~ sq ~ O    w    xq ~"sq ~sq ~sq ~$q ~ Qsq ~&q ~"sq ~sq ~$q ~ ?sq ~&q ~"sq ~+uq ~/   q ~"sq ~8sq ~<?@     q ~"q ~"xq ~"uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~"xq ~ Qq ~Wq ~E(�ysq ~Z�|�(   q ~aq ~jq ~iw   Csq ~Ȩ�sq ~ sq ~ sq ~ 
w   q ~pxq ~"q ~"sq ~ Eq ~ �sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~"sq ~sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~�q ~�uq ~>   q ~ Qq ~�q ~ ?q ~Wq ~ v��9�q ~�w   sq ~�O�sq ~ sq ~ sq ~ 
w   q ~pxq ~",q ~"+sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~"0sq ~sq ~sq ~$q ~ ?sq ~&q ~"3sq ~+uq ~/   q ~"3q ~"4q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �fv�sq ~ZȠU�   q ~aq ~eq ~iw   1sq ~@�m�sq ~ sq ~ sq ~ 
w   q ~zxq ~"<q ~";sq ~ Eq ~esq ~ L?z��    sq ~ sq ~ O   w   q ~ txq ~"@sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t?��q ~�w   Dsq ~��sq ~ sq ~ sq ~ 
w   q ~pq ~�xq ~"Nq ~"Msq ~ Eq ~�sq ~ Ll�    sq ~ sq ~ O   w   q ~ �q ~ ?xq ~"Rsq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?ڄs�q ~ew   6sq ~TB�|sq ~ sq ~ sq ~ 
w   q ~pxq ~"Zq ~"Ysq ~ Eq ~sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~"^sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?=�Pq ~ew   -sq ~�}]sq ~ sq ~ sq ~ 
w   q ~hxq ~"fq ~"esq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~"jsq ~sq ~sq ~$q ~ Qsq ~&q ~"msq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~"rsq ~+uq ~/   q ~"rsq ~8sq ~<?@     q ~"rq ~"mxq ~"muq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~"mxq ~ Qsq ~sq ~$q ~ ?sq ~&q ~"|sq ~+uq ~/   q ~"|q ~"}q ~�uq ~>   q ~ �q ~ `q ~Wq ~�q ~"yq ~huq ~>   q ~ Qq ~ �q ~ ?q ~Wq ~ vm���sq ~Z�ƥY   q ~eq ~jq ~iw   \sq ~b|�sq ~ sq ~ sq ~ 
w   q ~pxq ~"�q ~"�sq ~ Eq ~/sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~"�sq ~sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�sq ~8sq ~<?@     q ~�q ~�xq ~ ]uq ~>   q ~ `q ~ `q ~ Asq ~8sq ~<?@     q ~�xq ~ Qq ~Wq ~ t�]��q ~�w   sq ~I�Gmsq ~ sq ~ sq ~ 
w   q ~hxq ~"�q ~"�sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~"�sq ~sq ~sq ~$q ~ Qsq ~&q ~"�sq ~sq ~$q ~ �sq ~&q ~"�sq ~+uq ~/   sq ~sq ~$q ~ ?sq ~&q ~"�sq ~+uq ~/   q ~"�sq ~8sq ~<?@     q ~"�q ~"�xq ~"�uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~"�xq ~ Qsq ~sq ~$q ~ ?sq ~&q ~"�sq ~+uq ~/   q ~"�sq ~8sq ~<?@     q ~"�q ~"�xq ~"�uq ~>   q ~ ?q ~ ?sq ~8sq ~<?@     q ~"�xq ~ �sq ~8sq ~<?@     q ~"�q ~"�xq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~"�xq ~�q ~Wq ~��a��sq ~Z����   sq ~Z�ƥ�   q ~eq ~jq ~hq ~jq ~hw   Psq ~L�Zsq ~ sq ~ sq ~ 
w   q ~zq ~xq ~"�q ~"�sq ~ Eq ~sq ~ L�W9J    sq ~ sq ~ O   w   q ~ tq ~ �xq ~"�sq ~sq ~q ~Psq ~q ~Ssq ~+uq ~/   q ~aq ~dsq ~8sq ~<?@     q ~Pq ~Sxq ~zuq ~>   q ~ ?q ~ ?q ~ Asq ~8sq ~<?@     q ~Pxq ~ Qq ~Wq ~ tĊ��q ~bw   qsq ~�n9sq ~ sq ~ sq ~ 
w   q ~hq ~pxq ~"�q ~"�sq ~ Eq ~�sq ~ L�C�j    sq ~ sq ~ O   w   q ~�q ~ �xq ~"�sq ~sq ~q ~�sq ~q ~�sq ~q ~�sq ~+uq ~/   q ~�sq ~q ~�sq ~+uq ~/   q ~�q ~�q ~puq ~>   q ~ ?q ~ ?q ~Wq ~ �q ~�q ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~�xq ~ vq ~Wq ~Xsq ~8sq ~<?@      xq ~iw�Aq ~
w   zsq ~�CЭsq ~ sq ~ sq ~ 
w   q ~�xq ~"�q ~"�sq ~ Eq ~	#sq ~ L  E    sq ~ sq ~ O   w   q ~ ?xq ~"�sq ~wsq ~+uq ~/   q ~�q ~Wq ~ �uq ~>   q ~ �q ~ ;��Jq ~ew   Hsq ~W��sq ~ sq ~ sq ~ 
w   q ~pxq ~"�q ~"�sq ~ Eq ~�sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~"�sq ~wsq ~+uq ~/   q ~�q ~Wq ~puq ~>   q ~ ?q ~ ?�<�q ~ew   ;sq ~~��sq ~ sq ~ sq ~ 
w   q ~hxq ~#q ~#sq ~ Eq ~�sq ~ LW�m�    sq ~ sq ~ O   w   q ~�xq ~#	sq ~sq ~q ~sq ~q ~	sq ~q ~sq ~+uq ~/   q ~sq ~q ~sq ~+uq ~/   q ~q ~1q ~ fuq ~>   q ~ Qq ~ `sq ~8sq ~<?@     q ~q ~	xq ~�sq ~8sq ~<?@     q ~q ~	q ~xq ~huq ~>   q ~ Qq ~ �q ~ ?sq ~8sq ~<?@     q ~q ~	xq ~ vsq ~8sq ~<?@     q ~xq ~=q ~Wq ~?�8q ~Aw   psq ~�̱%sq ~ sq ~ sq ~ 
w   sq ~ 0q ~�t #0<e,<t,e>>t #0<e,<t,e>>:<e,<t,e>>xq ~# q ~#sq ~ Eq ~�sq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~#'sq ~sq ~sq ~$q ~ Qsq ~&q ~#*sq ~sq ~$q ~ ?sq ~&q ~#-sq ~+uq ~/   q ~#-sq ~+uq ~/   q ~#-sq ~8sq ~<?@     q ~#*q ~#-xq ~#*uq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~#*q ~#-xq ~#!uq ~>   q ~ ?q ~ Aq ~ ?sq ~8sq ~<?@     q ~#*xq ~ �q ~Wsq ~ 5JW'�t <<e,t>,<e,e>>q ~ Qq ~ ��K��sq ~Z��
�   q ~eq ~q ~iw   gsq ~/�sq ~ sq ~ sq ~ 
w   q ~pxq ~#Aq ~#@sq ~ Eq ~ �sq ~ L|!<    sq ~ sq ~ O   w   q ~ �xq ~#Esq ~wsq ~+uq ~/   q ~ �q ~Wq ~puq ~>   q ~ ?q ~ ?���q ~ew   +sq ~��Usq ~ sq ~ sq ~ 
w   q ~#!xq ~#Mq ~#Lsq ~ Eq ~	sq ~ L@M�4    sq ~ sq ~ O   w   q ~�xq ~#Qsq ~sq ~sq ~$q ~ Qsq ~&q ~#Tsq ~sq ~$q ~ ?sq ~&q ~#Wsq ~+uq ~/   q ~#Wsq ~+uq ~/   q ~#Wsq ~8sq ~<?@     q ~#Wq ~#Txq ~#Tuq ~>   q ~ ?q ~ Asq ~8sq ~<?@     q ~#Wq ~#Txq ~#!uq ~>   q ~ ?q ~ Aq ~ ?sq ~8sq ~<?@     q ~#Txq ~ �q ~Wq ~#;�N$!sq ~Z�7�   q ~esq ~ZȠU�   q ~aq ~eq ~hq ~iw   xsq ~ !        sr Yedu.cornell.cs.nlp.spf.parser.ccg.features.lambda.LogicalExpressionCoordinationFeatureSet�4tHWcg+ Z cpapFeaturesZ cpp1FeaturesZ reptFeaturesxpsr Dedu.cornell.cs.nlp.spf.parser.ccg.features.basic.RuleUsageFeatureSet�k�d�L2� D scaleZ unaryRulesOnlyL 	ignoreSetq ~ xp?������� sr java.util.HashSet�D�����4  xpw   ?@      xsr Ledu.cornell.cs.nlp.spf.parser.ccg.features.basic.DynamicWordSkippingFeatures%�q�� L emptyCategoryq ~L 
featureTagq ~ xpsq ~wp    sq ~`zT�lq ~bt EMPTYt DYNSKIPxq ~ sq ~ sq ~ O   w   q ~ xq ~#usr %java.util.Collections$UnmodifiableSet��я��U  xq ~ sq ~#lw   ?@     sr .edu.cornell.cs.nlp.spf.base.hashvector.KeyArgs���]e.ɘ I hashCodeL arg1q ~ L arg2q ~ L arg3q ~ L arg4q ~ L arg5q ~ xp2Iݬq ~ t 
TMPDEFAULTpppsq ~#ywzq ~ t XEMEDEFAULTpppsq ~#y'��q ~ t 
LEXDEFAULTpppxsr Bedu.cornell.cs.nlp.spf.ccg.lexicon.factored.lambda.FactoredLexicon�>�"z L lexemesq ~ (L lexemesByTypeq ~ (L 	templatesq ~ (xpsq ~ H?@     �w      zq ~msq ~#lw   ?@     q ~bq ~'q ~axq ~jsq ~#lw   ?@     q ~�q ~
q ~Rq ~�q ~	�q ~_q ~�q ~�q ~zq ~�q ~�xq ~�sq ~#lw   ?@     q ~�q ~q ~�xq ~�sq ~#lw   ?@     q ~|q ~
�q ~�xq ~.sq ~#lw   ?@     
q ~�q ~
�q ~�q ~�q ~q ~Dq ~<q ~�q ~�q ~#xq ~sq ~#lw   ?@     q ~xq ~<sq ~#lw   ?@     q ~1xq ~ sq ~#lw   ?@     q ~xq ~sq ~#lw    ?@     q ~�q ~�q ~�q ~q ~�q ~tq ~�q ~�q ~�q ~Uq ~�q ~�q ~�xq ~esq ~#lw   ?@     q ~Zq ~�q ~�q ~,q ~xq ~�xq ~>sq ~#lw   ?@     q ~3xq ~!sq ~#lw   ?@     q ~�q ~xq ~�sq ~#lw   ?@     q ~�q ~�q ~	xq ~
�sq ~#lw   ?@     q ~
|q ~3q ~xq ~�sq ~#lw   ?@     q ~�xq ~
sq ~#lw   ?@     q ~�q ~�q ~?xq ~sq ~#lw   ?@     q ~ xq ~�sq ~#lw   ?@     q ~�q ~�q ~_xq ~ xsq ~#lw   ?@     q ~,q ~Sq ~!q ~ Xq ~	lq ~�q ~�xq ~�sq ~#lw   ?@     q ~}xq ~�sq ~#lw   ?@     q ~�q ~xq ~	sq ~#lw   ?@     q ~	xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~�q ~zq ~�q ~xq ~
�sq ~#lw   ?@     q ~�q ~
�q ~[xq ~1sq ~#lw   ?@     q ~�q ~oq ~&xq ~�sq ~#lw    ?@     q ~�q ~�q ~xq ~�q ~$q ~�q ~ q ~+q ~�q ~�q ~�q ~]q ~�q ~�xq ~ �sq ~#lw   ?@     q ~�q ~dq ~ �xq ~�sq ~#lw   ?@     q ~Mq ~)q ~�xq ~sq ~#lw   ?@     q ~	q ~q ~xq ~sq ~#lw   ?@     q ~�q ~q ~	Vq ~�q ~	9xq ~)sq ~#lw   ?@     q ~xq ~<sq ~#lw   ?@     q ~�q ~�q ~1xq ~bsq ~#lw   ?@     q ~Tq ~�q ~xq ~=sq ~#lw   ?@     q ~ q ~�q ~3q ~�q ~	�q ~2q ~
Uq ~)q ~�q ~�q ~�q ~@xq ~0sq ~#lw   ?@     q ~q ~Sq ~%xq ~�sq ~#lw   ?@     q ~-q ~Oq ~�xq ~*sq ~#lw   ?@     q ~q ~�q ~wxq ~*sq ~#lw   ?@     q ~xq ~nsq ~#lw    ?@     q ~cq ~hq ~�q ~�q ~Dq ~�q ~�q ~�q ~'q ~�q ~Lq ~�q ~�q ~�xq ~�sq ~#lw   ?@     q ~�q ~5q ~�xq ~�sq ~#lw   ?@     q ~	�q ~	�q ~�xq ~'sq ~#lw   ?@     q ~q ~jq ~xq ~sq ~#lw   ?@     q ~�q ~�q ~ xq ~�sq ~#lw   ?@     q ~�q ~
-q ~�xq ~�sq ~#lw   ?@     q ~Sq ~�q ~q ~q ~xq ~<sq ~#lw   ?@     q ~�q ~ }q ~1xq ~sq ~#lw   ?@     q ~�xq ~_sq ~#lw   ?@     q ~�q ~$q ~Qxq ~�sq ~#lw   ?@     q ~�q ~�q ~�xq ~4sq ~#lw   ?@     q ~	Aq ~q ~)q ~�q ~wxq ~	�sq ~#lw   ?@     q ~aq ~	�q ~ �xq ~�sq ~#lw   ?@     q ~�q ~vq ~>xq ~sq ~#lw   ?@     q ~q ~	q ~,xq ~ Usq ~#lw   ?@     q ~xq ~�q ~Rq ~�q ~�q ~fq ~�q ~ +xq ~\sq ~#lw   ?@     q ~Qxq ~gsq ~#lw   ?@     q ~\xq ~sq ~#lw   ?@     q ~xq ~�sq ~#lw   ?@     q ~�q ~�q ~�xq ~$sq ~#lw   ?@     q ~�q ~
%q ~xq ~
sq ~#lw   ?@     q ~�q ~	�q ~�xq ~sq ~#lw   ?@     q ~�q ~xq ~Csq ~#lw   ?@     q ~�q ~
5q ~�q ~�q ~�q ~�q ~�q ~Bq ~Yq ~`q ~Sq ~4xq ~Psq ~#lw   ?@     q ~uq ~Eq ~pxq ~tsq ~#lw   ?@     q ~ixq ~�sq ~#lw   ?@     q ~�q ~�q ~�xq ~�sq ~#lw   ?@     q ~#q ~�q ~�xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~�xq ~	�sq ~#lw   ?@     q ~
�q ~Gq ~	�xq ~ �sq ~#lw   ?@     q ~�q ~ �q ~pxq ~�sq ~#lw    ?@     q ~}q ~q ~Yq ~�q ~mq ~�q ~�q ~
�q ~gq ~�q ~�q ~q ~
�q ~�q ~
Hq ~Bq ~4xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~�q ~�q ~ �q ~�q ~3q ~�q ~�xq ~sq ~#lw   ?@     q ~q ~�q ~9xq ~Vsq ~#lw   ?@     q ~Kxq ~	�sq ~#lw   ?@     q ~�q ~	�q ~�xq ~�sq ~#lw   ?@     q ~(q ~�q ~wxq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~�q ~�q ~�xq ~sq ~#lw   ?@     q ~
�q ~�xq ~�sq ~#lw   ?@     q ~	q ~�q ~�xq ~�sq ~#lw   ?@     q ~�q ~q ~sxq ~"sq ~#lw   ?@     q ~q ~q ~�xq ~Qsq ~#lw   ?@     q ~Cq ~�q ~�xq ~�sq ~#lw   ?@     q ~�xq ~:sq ~#lw   ?@     q ~/xq ~�sq ~#lw   ?@     q ~-q ~�q ~�xq ~�sq ~#lw   ?@     q ~Qq ~q ~�q ~Mxq ~Ksq ~#lw   ?@     q ~q ~@xq ~�sq ~#lw   ?@     q ~{xq ~�sq ~#lw   ?@     q ~�q ~�q ~
�xq ~�sq ~#lw   ?@     q ~	�q ~-q ~�xq ~xsq ~#lw   ?@     q ~�q ~jq ~�xq ~	�sq ~#lw   ?@     q ~	�q ~q ~xq ~�sq ~#lw   ?@     q ~�q ~`q ~�xq ~psq ~#lw   ?@     q ~�q ~eq ~�xq ~ �sq ~#lw   ?@     q ~ �q ~ �q ~
fxq ~jsq ~#lw   ?@     q ~�q ~Vq ~
�xq ~0sq ~#lw   ?@     q ~%xq ~sq ~#lw   ?@     q ~�xq ~|sq ~#lw   ?@     q ~qq ~�q ~axq ~	isq ~#lw   ?@     q ~�q ~gq ~	^xq ~
�sq ~#lw    ?@     q ~�q ~�q ~�q ~	�q ~Fq ~	Iq ~Bq ~q ~�q ~tq ~>q ~�q ~Fq ~q ~
�q ~cxq ~sq ~#lw   ?@     q ~�q ~q ~�xq ~#sq ~#lw   ?@     q ~oq ~q ~<xq ~sq ~#lw   ?@     q ~
�q ~�q ~ �xq ~'sq ~#lw   ?@     q ~8q ~q ~xq ~	6sq ~#lw   ?@     q ~	+xq ~
sq ~#lw    ?@     q ~�q ~>q ~Fq ~Bq ~cq ~

q ~�q ~8q ~Tq ~�q ~�q ~�q ~q ~jq ~xq ~	(sq ~#lw   ?@     q ~�q ~	q ~
xq ~sq ~#lw   ?@     q ~�q ~rq ~�xq ~Rsq ~#lw   ?@     q ~�q ~�q ~sq ~Eq ~�xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~
nq ~�xq ~sq ~#lw   ?@     q ~:q ~lq ~7q ~xq ~�sq ~#lw   ?@     q ~�q ~�q ~�q ~iq ~�q ~Oq ~Lxq ~	sq ~#lw   ?@     q ~lq ~�q ~	txq ~Psq ~#lw   ?@     q ~Eq ~�q ~�xq ~�sq ~#lw   ?@     q ~�q ~$q ~�xq ~�sq ~#lw   ?@     q ~wq ~�q ~[q ~�q ~�xq ~.sq ~#lw   ?@     q ~#xxsq ~ H?@     w       q ~sq ~#lw   ?@     q ~�q ~	q ~�q ~�q ~�xq ~ksq ~#lw   ?@     �q ~
�q ~-q ~�q ~�q ~�q ~�q ~q ~q ~�q ~�q ~�q ~
�q ~q ~�q ~
|q ~>q ~2q ~�q ~<q ~q ~Mq ~q ~�q ~mq ~#q ~ q ~	q ~ �q ~dq ~Yq ~�q ~
fq ~�q ~	q ~%q ~ �q ~�q ~�q ~�q ~�q ~sq ~�q ~�q ~�q ~gq ~�q ~�q ~)q ~q ~�q ~q ~	q ~�q ~4q ~�q ~>q ~�q ~Sq ~uq ~Bq ~q ~	�q ~
�q ~�q ~�q ~�q ~-q ~Uq ~�q ~	q ~�q ~�q ~�q ~	�q ~�q ~xq ~�q ~�q ~tq ~�q ~�q ~�q ~
�q ~cq ~�q ~Zq ~Fq ~q ~�q ~
Uq ~wq ~	tq ~cq ~'q ~�q ~ q ~�q ~	�q ~Qq ~eq ~�q ~q ~fq ~#q ~Yq ~�q ~�q ~�q ~�q ~%q ~�q ~wq ~jq ~1q ~	9q ~zq ~�q ~iq ~�q ~�q ~'q ~�q ~�q ~�q ~Oq ~�q ~
�q ~�q ~�q ~q ~:q ~
nq ~�q ~`q ~�q ~oq ~
-q ~�q ~xq ~	sq ~#lw   ?@     q ~�q ~�q ~wq ~�q ~�xq ~�sq ~#lw    ?@     q ~�q ~�q ~�q ~q ~�q ~\q ~�q ~/q ~q ~iq ~�q ~�q ~�q ~�q ~�q ~�q ~q ~ q ~�q ~}q ~�q ~	q ~3q ~Kxq ~�sq ~#lw   @?@     (q ~
�q ~8q ~�q ~	�q ~�q ~Qq ~pq ~�q ~_q ~�q ~�q ~oq ~Mq ~ �q ~lq ~q ~�q ~sq ~�q ~vq ~pq ~�q ~�q ~(q ~
%q ~�q ~�q ~	lq ~q ~�q ~�q ~q ~	�q ~�q ~�q ~Gq ~q ~�q ~�q ~xq ~ qsq ~#lw   ?@     q ~ Xxq ~ sq ~#lw   ?@     q ~�xq ~Xsq ~#lw   ?@     q ~Sxq ~Isq ~#lw   ?@     q ~	�q ~
�q ~Rq ~gq ~aq ~Dq ~q ~<q ~�q ~�q ~q ~axq ~�sq ~#lw   @?@     'q ~�q ~$q ~Eq ~q ~�q ~ �q ~
q ~�q ~ �q ~q ~Tq ~Sq ~q ~�q ~q ~�q ~q ~q ~Cq ~rq ~wq ~�q ~jq ~�q ~�q ~�q ~	�q ~)q ~�q ~[q ~�q ~�q ~�q ~�q ~>q ~�q ~
�q ~ �q ~xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   �?@     Wq ~�q ~�q ~	�q ~	�q ~�q ~lq ~�q ~Bq ~�q ~+q ~xq ~tq ~q ~[q ~�q ~
Hq ~7q ~Sq ~@q ~4q ~}q ~hq ~�q ~�q ~Bq ~ }q ~�q ~@q ~�q ~Vq ~qq ~�q ~�q ~�q ~�q ~Lq ~,q ~�q ~�q ~�q ~�q ~
�q ~Bq ~�q ~q ~�q ~�q ~5q ~�q ~xq ~3q ~q ~�q ~�q ~
�q ~q ~�q ~Tq ~�q ~�q ~�q ~cq ~�q ~�q ~�q ~�q ~3q ~Dq ~_q ~ �q ~�q ~	Iq ~Fq ~�q ~�q ~�q ~�q ~Qq ~q ~�q ~]q ~q ~Fq ~)q ~&q ~�q ~xq ~sq ~#lw   ?@     q ~q ~,q ~$q ~�q ~�q ~	+q ~�q ~xq ~ Msq ~#lw   ?@     q ~�q ~Rq ~3q ~ q ~�q ~ +xq ~	�sq ~#lw    ?@     q ~�q ~�q ~-q ~bq ~	�q ~�q ~	�q ~Eq ~q ~q ~�q ~,q ~q ~	^q ~�xq ~�sq ~#lw   ?@     q ~{xq ~&sq ~#lw   ?@     q ~!xq ~sq ~#lw   @?@     'q ~�q ~
5q ~�q ~�q ~�q ~�q ~�q ~Oq ~

q ~q ~1q ~8q ~Eq ~�q ~�q ~�q ~
�q ~�q ~Lq ~?q ~q ~�q ~zq ~�q ~$q ~�q ~�q ~�q ~|q ~�q ~�q ~�q ~�q ~�q ~�q ~`q ~�q ~jq ~9xq ~+sq ~#lw   ?@     q ~#q ~q ~1q ~axq ~�sq ~#lw   ?@     q ~q ~
q ~q ~�q ~�xq ~�sq ~#lw   ?@     q ~	Aq ~	Vq ~�q ~�q ~�xxsq ~ H?@     w       q ~!sq ~#lw   ?@     q ~!q ~�xq ~Msq ~#lw   �?@     3q ~ &q ~!�q ~�q ~#>q ~�q ~!q ~lq ~�q ~!�q ~�q ~�q ~�q ~"�q ~�q ~�q ~�q ~Hq ~�q ~q ~�q ~�q ~�q ~ Vq ~xq ~"Wq ~Fq ~ �q ~Tq ~�q ~")q ~�q ~*q ~�q ~!q ~"q ~�q ~Jq ~q ~ �q ~-q ~ 2q ~!Uq ~�q ~�q ~}q ~"�q ~<q ~�q ~Zq ~Dq ~�xq ~sq ~#lw   ?@     q ~�xq ~�sq ~#lw    ?@     q ~�q ~�q ~�q ~dq ~!�q ~ >q ~ �q ~�q ~�q ~-q ~q ~!�q ~�q ~�q ~lq ~"q ~�q ~ �q ~q ~cxq ~"�sq ~#lw   ?@     q ~�q ~�q ~!Bq ~"�xq ~ �sq ~#lw   ?@     q ~ �xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~�xq ~�sq ~#lw   ?@     q ~�q ~"�q ~�xq ~"Psq ~#lw   ?@     q ~"Kxq ~~sq ~#lw   ?@     q ~sxq ~�sq ~#lw    ?@     q ~q ~�q ~:q ~jq ~�q ~�q ~[q ~'q ~q ~�q ~"9q ~!-q ~�xq ~>sq ~#lw   ?@     q ~�q ~hq ~!aq ~q ~�q ~?q ~�q ~9xq ~@sq ~#lw   ?@     q ~8xq ~isq ~#lw    ?@     q ~"cq ~�q ~�q ~�q ~dq ~ bq ~#q ~"�q ~�q ~�q ~dq ~�q ~6xq ~^sq ~#lw   ?@     q ~Vxq ~Msq ~#lw   ?@     q ~Hxq ~#Osq ~#lw   ?@     q ~#q ~#Jxq ~�sq ~#lw   ?@     q ~ 
q ~�q ~�q ~Oxq ~�sq ~#lw   ?@     q ~�q ~�q ~q ~!�q ~"�q ~�q ~!�q ~�xq ~�sq ~#lw   ?@     q ~�xxsr 9edu.cornell.cs.nlp.spf.base.hashvector.FastTreeHashVector;��tQ57� L valuest 0Lit/unimi/dsi/fastutil/objects/Object2DoubleMap;xpsr 5it.unimi.dsi.fastutil.objects.Object2DoubleAVLTreeMap�7y�J| I countL storedComparatort Ljava/util/Comparator;xr <it.unimi.dsi.fastutil.objects.AbstractObject2DoubleSortedMap�c����  xr 6it.unimi.dsi.fastutil.objects.AbstractObject2DoubleMap�o��K<z  xr ;it.unimi.dsi.fastutil.objects.AbstractObject2DoubleFunction�o��K<z D defRetValuexp          Jpsq ~#yWD�t DYNSKIPppppw��      sq ~#yW�"�q ~ t LEXt 0t 0pw        sq ~#yW���q ~ q ~$5t 0t 35pw@$      sq ~#yW�&�q ~ q ~$5t 1t 1pw        sq ~#yW���q ~ q ~$5t 1t 13pw@$      sq ~#yW� �q ~ q ~$5t 10t 10pw        sq ~#yW�icq ~ q ~$5t 10t 3pw@$      sq ~#yW�i�q ~ q ~$5t 10t 8pw@$      sq ~#yZw,hq ~ q ~$5t 100t 11pw        sq ~#yZwC�q ~ q ~$5t 100t 78pw@5oz�G�sq ~#yZ�r�q ~ q ~$5t 101t 104pw@$      sq ~#yZ�sQq ~ q ~$5t 101t 107pw@$      sq ~#yZw8eq ~ q ~$5t 101t 37pw@$      sq ~#yZw?-q ~ q ~$5t 101t 51pw@$      sq ~#yZwC�q ~ q ~$5t 101t 67pw        sq ~#yZwJ�q ~ q ~$5t 101t 83pw@$      sq ~#yZwO)q ~ q ~$5t 101t 99pw@'���@nsq ~#yZw7�q ~ q ~$5t 102t 23pw        sq ~#yZw@%q ~ q ~$5t 102t 49pw@;�뤍sq ~#yZw?-q ~ q ~$5t 103t 31pw@$      sq ~#yZwC�q ~ q ~$5t 103t 48pw        sq ~#yZw<dq ~ q ~$5t 104t 19pw        sq ~#yZv�Tq ~ q ~$5t 104t 8pw@$      sq ~#yZw@q ~ q ~$5t 105t 18pw        sq ~#yZwC�q ~ q ~$5t 105t 27pw@$      sq ~#yZwV/q ~ q ~$5t 105t 75pw@$      sq ~#yZv�q ~ q ~$5t 105t 8pw?��s��֓sq ~#yZv�;q ~ q ~$5t 106t 3pw@5oz�G�sq ~#yZwRnq ~ q ~$5t 106t 55pw        sq ~#yZv��q ~ q ~$5t 106t 8pw@5oz�G�sq ~#yZwZMq ~ q ~$5t 107t 68pw        sq ~#yZwarq ~ q ~$5t 107t 85pw@$      sq ~#yZwRq ~ q ~$5t 108t 32pw        sq ~#yZwe3q ~ q ~$5t 108t 85pw@$      sq ~#yZ���q ~ q ~$5t 109t 137pw@$      sq ~#yZwa�q ~ q ~$5t 109t 69pw        sq ~#yZwd�q ~ q ~$5t 109t 72pw@$      sq ~#yW�$�q ~ q ~$5t 11t 11pw        sq ~#yW�?�q ~ q ~$5t 11t 87pw@5oz�G�sq ~#yZw�Bq ~ q ~$5t 110t 27pw@$      sq ~#yZv�3q ~ q ~$5t 110t 4pw        sq ~#yZw��q ~ q ~$5t 110t 75pw@$      sq ~#yZw�q ~ q ~$5t 111t 27pw@$      sq ~#yZw�q ~ q ~$5t 111t 55pw        sq ~#yZw��q ~ q ~$5t 111t 75pw@$      sq ~#yZw�Aq ~ q ~$5t 112t 19pw        sq ~#yZw��q ~ q ~$5t 112t 27pw@#��吢sq ~#yZw�Kq ~ q ~$5t 112t 75pw@$      sq ~#yZv�Wq ~ q ~$5t 113t 3pw@)I�L鼠sq ~#yZw��q ~ q ~$5t 113t 44pw        sq ~#yZw�Eq ~ q ~$5t 113t 49pw?�g�џ�sq ~#yZv��q ~ q ~$5t 113t 8pw@$      sq ~#yZw�Eq ~ q ~$5t 114t 39pw@$      sq ~#yZw�2q ~ q ~$5t 114t 70pw        sq ~#yZw�Lq ~ q ~$5t 115t 33pw        sq ~#yZw��q ~ q ~$5t 115t 81pw@$      sq ~#yZ���q ~ q ~$5t 116t 112pw@$      sq ~#yZw�-q ~ q ~$5t 116t 22pw@$      sq ~#yZw��q ~ q ~$5t 116t 71pw        sq ~#yZw�uq ~ q ~$5t 116t 80pw        sq ~#yZw�6q ~ q ~$5t 116t 90pw@$      sq ~#yZw¯q ~ q ~$5t 117t 32pw@$      sq ~#yZw��q ~ q ~$5t 117t 73pw        sq ~#yZw�Kq ~ q ~$5t 118t 15pw        sq ~#yZw�q ~ q ~$5t 118t 77pw@$      sq ~#yZw:q ~ q ~$5t 119t 6pw@$      sq ~#yW�(�q ~ q ~$5t 12t 12pw        sq ~#yW�)Rq ~ q ~$5t 12t 17pw        sq ~#yW�8Vq ~ q ~$5t 12t 57pw@$      sq ~#yZx�q ~ q ~$5t 120t 17pw@$      sq ~#yZx �q ~ q ~$5t 120t 44pw@$      sq ~#yZx!aq ~ q ~$5t 120t 49pw        sq ~#yZ�[�q ~ q ~$5t 121t 106pw        sq ~#yZ�\q ~ q ~$5t 121t 107pw        sq ~#yZx/�q ~ q ~$5t 121t 74pw        sq ~#yZx3lq ~ q ~$5t 121t 83pw@$      sq ~#yZx7�q ~ q ~$5t 121t 98pw@$      sq ~#yZx7�q ~ q ~$5t 121t 99pw@'���@nsq ~#yZx!#q ~ q ~$5t 122t 27pw@$      sq ~#yZx%"q ~ q ~$5t 122t 39pw        sq ~#yZx3�q ~ q ~$5t 122t 75pw@$      sq ~#yZwhxq ~ q ~$5t 123t 1pw        sq ~#yZx$�q ~ q ~$5t 123t 27pw@"
\�Hq�sq ~#yZx7kq ~ q ~$5t 123t 75pw@$      sq ~#yZ�f�q ~ q ~$5t 124t 102pw        sq ~#yZ�jYq ~ q ~$5t 124t 111pw@$      sq ~#yZx(
q ~ q ~$5t 124t 22pw@$      sq ~#yZx7Lq ~ q ~$5t 124t 64pw@$      sq ~#yZx;Kq ~ q ~$5t 124t 76pw        sq ~#yZxB�q ~ q ~$5t 124t 97pw@$      sq ~#yZwp8q ~ q ~$5t 125t 3pw@$      sq ~#yZx/�q ~ q ~$5t 125t 35pw        sq ~#yZwp�q ~ q ~$5t 125t 8pw@$      sq ~#yZws�q ~ q ~$5t 126t 0pw@%U�i�g�sq ~#yZxB�q ~ q ~$5t 126t 75pw        sq ~#yZx/�q ~ q ~$5t 127t 15pw        sq ~#yZx0q ~ q ~$5t 127t 16pw@$      sq ~#yZw{{q ~ q ~$5t 128t 3pw@$      sq ~#yZx;q ~ q ~$5t 128t 34pw        sq ~#yZw|q ~ q ~$5t 128t 8pw@$      sq ~#yZxI�q ~ q ~$5t 129t 60pw        sq ~#yZxQ�q ~ q ~$5t 129t 85pw@$      sq ~#yW�,�q ~ q ~$5t 13t 13pw        sq ~#yW�;�q ~ q ~$5t 13t 55pw@$      sq ~#yZx�cq ~ q ~$5t 130t 46pw@$      sq ~#yZx�Cq ~ q ~$5t 130t 57pw        sq ~#yZx��q ~ q ~$5t 131t 60pw        sq ~#yZw�q ~ q ~$5t 131t 7pw@$      sq ~#yZw��q ~ q ~$5t 132t 7pw        sq ~#yZx��q ~ q ~$5t 132t 85pw@$      sq ~#yZ��3q ~ q ~$5t 133t 137pw@5oz�G�sq ~#yZx��q ~ q ~$5t 133t 69pw@5oz�G�sq ~#yZx�Fq ~ q ~$5t 133t 79pw        sq ~#yZx��q ~ q ~$5t 134t 38pw@$      sq ~#yZw�3q ~ q ~$5t 134t 6pw        sq ~#yZx��q ~ q ~$5t 135t 27pw@#]<6(��sq ~#yZx��q ~ q ~$5t 135t 66pw        sq ~#yZx�Lq ~ q ~$5t 135t 75pw@$      sq ~#yZw�Xq ~ q ~$5t 136t 3pw@5oz�G�sq ~#yZx�q ~ q ~$5t 136t 75pw        sq ~#yZw��q ~ q ~$5t 136t 8pw@5oz�G�sq ~#yZ��xq ~ q ~$5t 137t 103pw@$      sq ~#yZw�Wq ~ q ~$5t 137t 5pw@$      sq ~#yZx��q ~ q ~$5t 138t 19pw        sq ~#yZx�q ~ q ~$5t 138t 27pw@$      sq ~#yZx��q ~ q ~$5t 138t 75pw@$      sq ~#yZx�Mq ~ q ~$5t 139t 23pw        sq ~#yZx��q ~ q ~$5t 139t 27pw@$      sq ~#yZx�Pq ~ q ~$5t 139t 75pw@$      sq ~#yW�0wq ~ q ~$5t 14t 14pw        sq ~#yW�7�q ~ q ~$5t 14t 32pw@$      sq ~#yZy�q ~ q ~$5t 140t 61pw        sq ~#yZy�q ~ q ~$5t 140t 85pw@$      sq ~#yZy�q ~ q ~$5t 140t 86pw@$      sq ~#yZxI�q ~ q ~$5t 141t 2pw        sq ~#yZxJq ~ q ~$5t 141t 4pw@$      sq ~#yZ�S�q ~ q ~$5t 142t 137pw@$      sq ~#yZy#q ~ q ~$5t 142t 69pw        sq ~#yZyq ~ q ~$5t 142t 72pw@$      sq ~#yZy�q ~ q ~$5t 143t 27pw@$      sq ~#yZy�q ~ q ~$5t 143t 39pw        sq ~#yZy )q ~ q ~$5t 143t 75pw@$      sq ~#yZxU5q ~ q ~$5t 144t 3pw@$      sq ~#yZy+q ~ q ~$5t 144t 41pw        sq ~#yZxU�q ~ q ~$5t 144t 8pw@$      sq ~#yZy'mq ~ q ~$5t 145t 73pw@$      sq ~#yZx\�q ~ q ~$5t 146t 3pw@$      sq ~#yZx\�q ~ q ~$5t 146t 4pw        sq ~#yZx]Rq ~ q ~$5t 146t 8pw@$      sq ~#yZ�f�q ~ q ~$5t 147t 137pw@$�)�o�Usq ~#yZy+�q ~ q ~$5t 147t 69pw@(�5&h�hsq ~#yZy/�q ~ q ~$5t 147t 79pw        sq ~#yZy*�q ~ q ~$5t 148t 50pw        sq ~#yZxd�q ~ q ~$5t 148t 8pw@$      sq ~#yZy gq ~ q ~$5t 149t 17pw        sq ~#yZy �q ~ q ~$5t 149t 19pw@$      sq ~#yZy+q ~ q ~$5t 149t 42pw@$      sq ~#yZy.�q ~ q ~$5t 149t 52pw@$      sq ~#yW�4vq ~ q ~$5t 15t 16pw        sq ~#yW�|(q ~ q ~$5t 15t 3pw@$      sq ~#yW�;]q ~ q ~$5t 15t 31pw        sq ~#yW�|�q ~ q ~$5t 15t 8pw@$      sq ~#yZx�+q ~ q ~$5t 150t 8pw@$      sq ~#yZy��q ~ q ~$5t 150t 81pw        sq ~#yZy}�q ~ q ~$5t 151t 34pw        sq ~#yZx��q ~ q ~$5t 151t 8pw@$      sq ~#yZy�Jq ~ q ~$5t 152t 83pw@$      sq ~#yZy��q ~ q ~$5t 152t 98pw        sq ~#yZy��q ~ q ~$5t 152t 99pw@(1���ssq ~#yZ���q ~ q ~$5t 153t 137pw@$      sq ~#yZy�+q ~ q ~$5t 153t 72pw@$      sq ~#yZy�q ~ q ~$5t 153t 79pw        sq ~#yZy��q ~ q ~$5t 154t 26pw@!��Hsq ~#yZy�cq ~ q ~$5t 154t 48pw        sq ~#yZy��q ~ q ~$5t 154t 66pw@/��!'sq ~#yZy��q ~ q ~$5t 155t 18pw        sq ~#yZx��q ~ q ~$5t 155t 8pw@$      sq ~#yZy�*q ~ q ~$5t 156t 54pw@$      sq ~#yZx�zq ~ q ~$5t 157t 0pw        sq ~#yZx��q ~ q ~$5t 157t 3pw@$      sq ~#yZx�rq ~ q ~$5t 157t 8pw@$      sq ~#yZ���q ~ q ~$5t 158t 115pw        sq ~#yZy��q ~ q ~$5t 158t 84pw@5oz�G�sq ~#yZy��q ~ q ~$5t 159t 17pw        sq ~#yZx�Yq ~ q ~$5t 159t 3pw@$      sq ~#yZx��q ~ q ~$5t 159t 8pw@$      sq ~#yW�7�q ~ q ~$5t 16t 14pw        sq ~#yW�Gyq ~ q ~$5t 16t 58pw@$      sq ~#yZy.�q ~ q ~$5t 160t 3pw@$      sq ~#yZy�"q ~ q ~$5t 160t 55pw        sq ~#yZy/�q ~ q ~$5t 160t 8pw@$      sq ~#yZ�-�q ~ q ~$5t 161t 107pw@��ыsq ~#yZy�q ~ q ~$5t 161t 37pw        sq ~#yZzFq ~ q ~$5t 161t 74pw@$      sq ~#yZy�q ~ q ~$5t 162t 58pw��3H4�rjsq ~#yZz�q ~ q ~$5t 162t 73pw@$      sq ~#yZz�q ~ q ~$5t 162t 85pw@�Xx'sq ~#yZz	q ~ q ~$5t 162t 86pw        sq ~#yZy:�q ~ q ~$5t 163t 7pw@$      sq ~#yZz�q ~ q ~$5t 163t 85pw        sq ~#yZzjq ~ q ~$5t 164t 73pw        sq ~#yZziq ~ q ~$5t 164t 85pw@$      sq ~#yZz�q ~ q ~$5t 164t 86pw@$      sq ~#yZzhq ~ q ~$5t 165t 87pw        sq ~#yZz�q ~ q ~$5t 165t 93pw@%��9�}qsq ~#yZyEuq ~ q ~$5t 166t 3pw@$      sq ~#yZz�q ~ q ~$5t 166t 66pw        sq ~#yZyFq ~ q ~$5t 166t 8pw@$      sq ~#yZzeq ~ q ~$5t 167t 15pw        sq ~#yZzdq ~ q ~$5t 167t 27pw@&eNO���sq ~#yZz�q ~ q ~$5t 167t 75pw@$      sq ~#yZz	q ~ q ~$5t 168t 26pw@&Q��/(sq ~#yZziq ~ q ~$5t 168t 45pw        sq ~#yZz+q ~ q ~$5t 169t 33pw@$      sq ~#yZz�q ~ q ~$5t 169t 40pw        sq ~#yW�<6q ~ q ~$5t 17t 18pw        sq ~#yWă�q ~ q ~$5t 17t 3pw@$      sq ~#yWĄEq ~ q ~$5t 17t 8pw@$      sq ~#yZzc{q ~ q ~$5t 170t 39pw        sq ~#yZzfcq ~ q ~$5t 170t 42pw@$      sq ~#yZzn�q ~ q ~$5t 171t 59pw        sq ~#yZy��q ~ q ~$5t 171t 8pw@$      sq ~#yZ���q ~ q ~$5t 172t 119pw@5oz�G�sq ~#yZ��Tq ~ q ~$5t 172t 120pw@5oz�G�sq ~#yZz}�q ~ q ~$5t 172t 88pw        sq ~#yZy��q ~ q ~$5t 173t 3pw@$      sq ~#yZzv@q ~ q ~$5t 173t 59pw        sq ~#yZy�,q ~ q ~$5t 173t 8pw@$      sq ~#yZzyfq ~ q ~$5t 174t 54pw@$      sq ~#yZzrAq ~ q ~$5t 175t 27pw��N>)L�&sq ~#yZzy(q ~ q ~$5t 175t 42pw@�e��'�sq ~#yZz�&q ~ q ~$5t 175t 66pw        sq ~#yZzu�q ~ q ~$5t 176t 24pw@$      sq ~#yZzy�q ~ q ~$5t 176t 35pw        sq ~#yZz|�q ~ q ~$5t 177t 32pw@$      sq ~#yZy�Oq ~ q ~$5t 177t 9pw        sq ~#yZzx�q ~ q ~$5t 178t 10pw@$      sq ~#yZy�Vq ~ q ~$5t 178t 3pw        sq ~#yZz�Lq ~ q ~$5t 178t 41pw@$      sq ~#yZz�kq ~ q ~$5t 179t 32pw        sq ~#yZz��q ~ q ~$5t 179t 85pw@$      sq ~#yW�@q ~ q ~$5t 18t 19pw        sq ~#yW�K:q ~ q ~$5t 18t 48pw@$      sq ~#yZz�}q ~ q ~$5t 180t 36pw        sq ~#yZz�#q ~ q ~$5t 180t 85pw@$      sq ~#yZz�q ~ q ~$5t 181t 7pw        sq ~#yZz��q ~ q ~$5t 181t 73pw@$      sq ~#yZ��q ~ q ~$5t 182t 103pw@$      sq ~#yZzmq ~ q ~$5t 182t 5pw@$      sq ~#yZzރq ~ q ~$5t 183t 22pw@$      sq ~#yZz��q ~ q ~$5t 183t 89pw        sq ~#yZ�!�q ~ q ~$5t 184t 109pw@5oz�G�sq ~#yZz�q ~ q ~$5t 184t 37pw        sq ~#yZ{ -q ~ q ~$5t 185t 91pw@$      sq ~#yZz�aq ~ q ~$5t 186t 27pw@$      sq ~#yZz�Hq ~ q ~$5t 186t 42pw        sq ~#yZz��q ~ q ~$5t 186t 75pw@$      sq ~#yZ{jq ~ q ~$5t 187t 85pw@$      sq ~#yZ{�q ~ q ~$5t 187t 86pw@$      sq ~#yZ�0qq ~ q ~$5t 188t 106pw@$      sq ~#yZ�0�q ~ q ~$5t 188t 109pw@$      sq ~#yZ{�q ~ q ~$5t 188t 78pw@$      sq ~#yZ�?�q ~ q ~$5t 189t 137pw@$      sq ~#yZ{�q ~ q ~$5t 189t 72pw@$      sq ~#yZ{�q ~ q ~$5t 189t 79pw        sq ~#yW�F�q ~ q ~$5t 19t 20pw        sq ~#yWċ,q ~ q ~$5t 19t 3pw@$      sq ~#yWċ�q ~ q ~$5t 19t 8pw@%��9�}qsq ~#yZ{L9q ~ q ~$5t 190t 39pw        sq ~#yZz��q ~ q ~$5t 190t 8pw@5v��n�sq ~#yZz�Iq ~ q ~$5t 191t 7pw        sq ~#yZ{bCq ~ q ~$5t 191t 85pw@5oz�G�sq ~#yZ��oq ~ q ~$5t 192t 123pw@$      sq ~#yZ{i�q ~ q ~$5t 192t 94pw@$      sq ~#yZ{b�q ~ q ~$5t 193t 67pw@$      sq ~#yZ{Z�q ~ q ~$5t 194t 36pw        sq ~#yZ{m�q ~ q ~$5t 194t 85pw@$      sq ~#yZ{m�q ~ q ~$5t 194t 86pw@$      sq ~#yZ{ZEq ~ q ~$5t 195t 21pw        sq ~#yZ{qGq ~ q ~$5t 195t 85pw@$      sq ~#yZ���q ~ q ~$5t 196t 130pw@5oz�G�sq ~#yZ{x�q ~ q ~$5t 196t 95pw@5oz�G�sq ~#yZ{y&q ~ q ~$5t 197t 88pw@@�鹙�sq ~#yZ{|�q ~ q ~$5t 197t 96pw        sq ~#yZ{|�q ~ q ~$5t 198t 85pw@$      sq ~#yZ{faq ~ q ~$5t 199t 18pw        sq ~#yZz��q ~ q ~$5t 199t 3pw@$      sq ~#yZz�pq ~ q ~$5t 199t 8pw@$      sq ~#yW�*�q ~ q ~$5t 2t 2pw        sq ~#yW��lq ~ q ~$5t 2t 63pw@$      sq ~#yWř6q ~ q ~$5t 20t 21pw        sq ~#yWŝ�q ~ q ~$5t 20t 36pw        sq ~#yWŰ8q ~ q ~$5t 20t 85pw@5oz�G�sq ~#yZ�Z�q ~ q ~$5t 200t 73pw        sq ~#yZ�^�q ~ q ~$5t 200t 85pw@@�鹙�sq ~#yZ�L%q ~ q ~$5t 201t 27pw@$      sq ~#yZ�O,q ~ q ~$5t 201t 31pw        sq ~#yZ�^�q ~ q ~$5t 201t 75pw@$      sq ~#yZ���q ~ q ~$5t 202t 109pw@5oz�G�sq ~#yZ�S�q ~ q ~$5t 202t 37pw        sq ~#yZ�Sq ~ q ~$5t 203t 22pw@$      sq ~#yZ�bNq ~ q ~$5t 203t 64pw        sq ~#yZ�R�q ~ q ~$5t 204t 11pw@$      sq ~#yZ�e�q ~ q ~$5t 204t 62pw@$      sq ~#yZ�q3q ~ q ~$5t 204t 93pw@'���@nsq ~#yZ�mrq ~ q ~$5t 205t 73pw        sq ~#yZ�qqq ~ q ~$5t 205t 85pw@$      sq ~#yZ�u2q ~ q ~$5t 206t 85pw@$      sq ~#yZ�uQq ~ q ~$5t 206t 86pw@$      sq ~#yZ�p�q ~ q ~$5t 207t 61pw        sq ~#yZ�x�q ~ q ~$5t 207t 85pw@$      sq ~#yZ��_q ~ q ~$5t 208t 101pw        sq ~#yZ�f�q ~ q ~$5t 208t 29pw        sq ~#yZ�|vq ~ q ~$5t 208t 83pw@$      sq ~#yZ���q ~ q ~$5t 209t 119pw        sq ~#yZ���q ~ q ~$5t 209t 121pw@5oz�G�sq ~#yZ���q ~ q ~$5t 209t 129pw@5oz�G�sq ~#yZ��Uq ~ q ~$5t 209t 96pw        sq ~#yW���q ~ q ~$5t 21t 102pw@$      sq ~#yWŝq ~ q ~$5t 21t 22pw@$      sq ~#yWů�q ~ q ~$5t 21t 71pw@$      sq ~#yWŰWq ~ q ~$5t 21t 76pw@$      sq ~#yWŷ]q ~ q ~$5t 21t 92pw        sq ~#yZ��	q ~ q ~$5t 210t 21pw        sq ~#yZ��q ~ q ~$5t 210t 85pw@$      sq ~#yZ��*q ~ q ~$5t 210t 86pw@$      sq ~#yZ���q ~ q ~$5t 211t 18pw@$      sq ~#yZ���q ~ q ~$5t 211t 20pw        sq ~#yZ��Eq ~ q ~$5t 212t 27pw@$      sq ~#yZ��jq ~ q ~$5t 212t 44pw        sq ~#yZ���q ~ q ~$5t 212t 75pw@$      sq ~#yZ��Dq ~ q ~$5t 213t 29pw        sq ~#yZ�ҏq ~ q ~$5t 213t 51pw@$      sq ~#yZ��q ~ q ~$5t 214t 3pw@$      sq ~#yZ���q ~ q ~$5t 214t 44pw        sq ~#yZ�4q ~ q ~$5t 214t 8pw@$      sq ~#yZ���q ~ q ~$5t 215t 73pw        sq ~#yZ���q ~ q ~$5t 215t 85pw@5oz�G�sq ~#yZ�9q ~ q ~$5t 216t 137pw@$      sq ~#yZ��q ~ q ~$5t 216t 69pw@$      sq ~#yZ� �q ~ q ~$5t 217t 137pw@$      sq ~#yZ��4q ~ q ~$5t 217t 72pw@$      sq ~#yZ��q ~ q ~$5t 217t 79pw        sq ~#yZ�q ~ q ~$5t 218t 111pw@$      sq ~#yZ��q ~ q ~$5t 218t 112pw        sq ~#yZ�q ~ q ~$5t 218t 116pw        sq ~#yZ��0q ~ q ~$5t 218t 22pw@$      sq ~#yZ��q ~ q ~$5t 218t 89pw@$      sq ~#yZ��wq ~ q ~$5t 218t 92pw        sq ~#yZ��Nq ~ q ~$5t 219t 25pw        sq ~#yZ�"�q ~ q ~$5t 219t 8pw@$      sq ~#yWŠ�q ~ q ~$5t 22t 23pw        sq ~#yWŨq ~ q ~$5t 22t 40pw@$      sq ~#yZ�<�q ~ q ~$5t 220t 58pw        sq ~#yZ�Gjq ~ q ~$5t 220t 85pw@$      sq ~#yZ�G�q ~ q ~$5t 220t 86pw@$      sq ~#yZ�0�q ~ q ~$5t 221t 14pw        sq ~#yZ�K+q ~ q ~$5t 221t 85pw@$      sq ~#yZ�4�q ~ q ~$5t 222t 14pw        sq ~#yZ�F�q ~ q ~$5t 222t 60pw@$      sq ~#yZ�R�q ~ q ~$5t 223t 85pw@5oz�G�sq ~#yZ���q ~ q ~$5t 223t 9pw        sq ~#yZ�Vnq ~ q ~$5t 224t 85pw@$      sq ~#yZ��q ~ q ~$5t 225t 103pw@$      sq ~#yZ���q ~ q ~$5t 225t 5pw@$      sq ~#yZ�J�q ~ q ~$5t 226t 32pw@$      sq ~#yZ�Y�q ~ q ~$5t 226t 73pw        sq ~#yZ��;q ~ q ~$5t 227t 3pw@5oz�G�sq ~#yZ�Npq ~ q ~$5t 227t 31pw        sq ~#yZ���q ~ q ~$5t 227t 8pw@5oz�G�sq ~#yZ�Zq ~ q ~$5t 228t 54pw@%Sx�d��sq ~#yZ���q ~ q ~$5t 229t 2pw        sq ~#yZ���q ~ q ~$5t 229t 3pw@$      sq ~#yZ��Xq ~ q ~$5t 229t 8pw@$      sq ~#yWŠ�q ~ q ~$5t 23t 12pw@$      sq ~#yWŤ�q ~ q ~$5t 23t 24pw        sq ~#yWŬ�q ~ q ~$5t 23t 47pw        sq ~#yZ��q ~ q ~$5t 230t 103pw@$      sq ~#yZ��q ~ q ~$5t 230t 5pw@$      sq ~#yZ��q ~ q ~$5t 231t 104pw        sq ~#yZ���q ~ q ~$5t 231t 107pw@$      sq ~#yZ���q ~ q ~$5t 232t 25pw        sq ~#yZ���q ~ q ~$5t 232t 47pw@$      sq ~#yZ��q ~ q ~$5t 233t 85pw@$      sq ~#yZ��+q ~ q ~$5t 233t 86pw@$      sq ~#yZ���q ~ q ~$5t 234t 27pw@$      sq ~#yZ���q ~ q ~$5t 234t 6pw        sq ~#yZ��q ~ q ~$5t 234t 75pw@$      sq ~#yZ�6q ~ q ~$5t 235t 137pw@$      sq ~#yZ�ǈq ~ q ~$5t 235t 69pw        sq ~#yZ��pq ~ q ~$5t 235t 72pw@$      sq ~#yZ��vq ~ q ~$5t 236t 105pw@$      sq ~#yZ��q ~ q ~$5t 237t 85pw@$      sq ~#yZ�Tq ~ q ~$5t 237t 9pw        sq ~#yZ�Ҭq ~ q ~$5t 238t 68pw        sq ~#yZ�q ~ q ~$5t 238t 9pw@5oz�G�sq ~#yZ�:q ~ q ~$5t 239t 137pw@5oz�G�sq ~#yZ�֌q ~ q ~$5t 239t 69pw@5oz�G�sq ~#yWũq ~ q ~$5t 24t 28pw        sq ~#yW���q ~ q ~$5t 24t 4pw        sq ~#yWŷ�q ~ q ~$5t 24t 66pw@F�U�i�sq ~#yZ�[�q ~ q ~$5t 240t 112pw@5oz�G�sq ~#yZ�0�q ~ q ~$5t 240t 89pw        sq ~#yZ�3Nq ~ q ~$5t 240t 90pw@5oz�G�sq ~#yZ�)q ~ q ~$5t 241t 58pw        sq ~#yZ�3�q ~ q ~$5t 241t 85pw@$      sq ~#yZ�4q ~ q ~$5t 241t 86pw@$      sq ~#yZ�/�q ~ q ~$5t 242t 60pw@$      sq ~#yZ�7�q ~ q ~$5t 242t 85pw        sq ~#yZ�0�q ~ q ~$5t 243t 58pw        sq ~#yZ�;kq ~ q ~$5t 243t 85pw@$      sq ~#yZ�;�q ~ q ~$5t 243t 86pw@$      sq ~#yZ�g�q ~ q ~$5t 244t 108pw@@�鹙�sq ~#yZ�jyq ~ q ~$5t 245t 100pw@$      sq ~#yZ�k�q ~ q ~$5t 245t 109pw        sq ~#yZ�C+q ~ q ~$5t 245t 87pw@$      sq ~#yZ�7Mq ~ q ~$5t 246t 42pw@$      sq ~#yZ�BRq ~ q ~$5t 246t 70pw        sq ~#yZ�~q ~ q ~$5t 247t 137pw@$      sq ~#yZ�Ciq ~ q ~$5t 247t 69pw        sq ~#yZ�FQq ~ q ~$5t 247t 72pw@%U��kK�sq ~#yZ�y}q ~ q ~$5t 248t 110pw@$      sq ~#yZ�U6q ~ q ~$5t 249t 91pw@$      sq ~#yWŨ�q ~ q ~$5t 25t 17pw        sq ~#yWŬ�q ~ q ~$5t 25t 27pw@$      sq ~#yWſ<q ~ q ~$5t 25t 75pw@$      sq ~#yZ���q ~ q ~$5t 250t 36pw@@�鹙�sq ~#yZ���q ~ q ~$5t 250t 58pw        sq ~#yZ��1q ~ q ~$5t 251t 103pw@5oz�G�sq ~#yZ��q ~ q ~$5t 251t 5pw@5oz�G�sq ~#yZ��#q ~ q ~$5t 252t 58pw        sq ~#yZ���q ~ q ~$5t 252t 60pw@$      sq ~#yZ��rq ~ q ~$5t 253t 137pw@5oz�G�sq ~#yZ���q ~ q ~$5t 253t 69pw@5oz�G�sq ~#yZ���q ~ q ~$5t 253t 72pw        sq ~#yZ���q ~ q ~$5t 254t 111pw@$      sq ~#yZ�ߒq ~ q ~$5t 254t 116pw@$      sq ~#yZ���q ~ q ~$5t 254t 22pw@$      sq ~#yZ��Nq ~ q ~$5t 254t 71pw@!��B��sq ~#yZ���q ~ q ~$5t 254t 76pw@$      sq ~#yZ���q ~ q ~$5t 254t 92pw@!��B��sq ~#yZ���q ~ q ~$5t 254t 97pw@!��B��sq ~#yZ��Jq ~ q ~$5t 255t 21pw@$      sq ~#yZ��*q ~ q ~$5t 255t 32pw        sq ~#yZ��Nq ~ q ~$5t 255t 61pw@$      sq ~#yZ��'q ~ q ~$5t 255t 68pw@$      sq ~#yZ��'q ~ q ~$5t 256t 58pw        sq ~#yZ��q ~ q ~$5t 256t 85pw@$      sq ~#yZ���q ~ q ~$5t 257t 73pw@$      sq ~#yZ��q ~ q ~$5t 257t 9pw        sq ~#yZ���q ~ q ~$5t 258t 22pw@$      sq ~#yZ���q ~ q ~$5t 258t 64pw@$      sq ~#yZ��9q ~ q ~$5t 259t 103pw@@�鹙�sq ~#yZ��q ~ q ~$5t 259t 5pw@@�鹙�sq ~#yWŬ�q ~ q ~$5t 26t 16pw        sq ~#yW��Hq ~ q ~$5t 26t 3pw@$      sq ~#yW���q ~ q ~$5t 26t 8pw@$      sq ~#yZ�L�q ~ q ~$5t 260t 137pw@$      sq ~#yZ��q ~ q ~$5t 260t 69pw@ �Q,4�sq ~#yZ��q ~ q ~$5t 260t 72pw        sq ~#yZ��q ~ q ~$5t 261t 72pw        sq ~#yZ�bq ~ q ~$5t 261t 79pw@@�鹙�sq ~#yZ�O�q ~ q ~$5t 262t 124pw@i���sq ~#yZ��q ~ q ~$5t 262t 65pw        sq ~#yZ�Lq ~ q ~$5t 263t 103pw@$      sq ~#yZ�Q�q ~ q ~$5t 263t 5pw@$      sq ~#yZ� �q ~ q ~$5t 264t 69pw        sq ~#yZ�#�q ~ q ~$5t 264t 72pw@@�鹙�sq ~#yZ� Iq ~ q ~$5t 265t 54pw@$      sq ~#yZ�/lq ~ q ~$5t 266t 85pw@5oz�G�sq ~#yZ�^�q ~ q ~$5t 267t 113pw@5oz�G�sq ~#yZ�_Sq ~ q ~$5t 267t 117pw        sq ~#yZ�fq ~ q ~$5t 267t 131pw@5oz�G�sq ~#yZ�byq ~ q ~$5t 268t 112pw@5oz�G�sq ~#yZ�:q ~ q ~$5t 268t 90pw@5oz�G�sq ~#yZ�2�q ~ q ~$5t 269t 60pw        sq ~#yZ�:�q ~ q ~$5t 269t 85pw@$      sq ~#yZ�:�q ~ q ~$5t 269t 86pw@$      sq ~#yWų�q ~ q ~$5t 27t 25pw        sq ~#yW��	q ~ q ~$5t 27t 3pw@$o� �@�sq ~#yWſ�q ~ q ~$5t 27t 59pw        sq ~#yW���q ~ q ~$5t 27t 8pw@$      sq ~#yZ��-q ~ q ~$5t 270t 115pw@$      sq ~#yZ���q ~ q ~$5t 270t 94pw        sq ~#yZ�Įq ~ q ~$5t 271t 137pw@$      sq ~#yZ�� q ~ q ~$5t 271t 69pw        sq ~#yZ���q ~ q ~$5t 271t 72pw@$      sq ~#yZ�}�q ~ q ~$5t 272t 22pw@$      sq ~#yZ��&q ~ q ~$5t 272t 64pw��Oy���sq ~#yZ���q ~ q ~$5t 272t 71pw���&��N�sq ~#yZ��Cq ~ q ~$5t 272t 89pw��Oy���sq ~#yZ��+q ~ q ~$5t 272t 92pw���&��N�sq ~#yZ���q ~ q ~$5t 272t 97pw���&��N�sq ~#yZ��Qq ~ q ~$5t 273t 114pw@$      sq ~#yZ�Įq ~ q ~$5t 273t 117pw@$      sq ~#yZ��vq ~ q ~$5t 273t 131pw        sq ~#yZ��'q ~ q ~$5t 274t 32pw@$      sq ~#yZ���q ~ q ~$5t 274t 36pw        sq ~#yZ�Ӳq ~ q ~$5t 275t 137pw@$      sq ~#yZ���q ~ q ~$5t 275t 72pw@$      sq ~#yZ���q ~ q ~$5t 275t 79pw        sq ~#yZ���q ~ q ~$5t 276t 73pw        sq ~#yZ���q ~ q ~$5t 276t 85pw@$      sq ~#yZ���q ~ q ~$5t 276t 86pw@$      sq ~#yZ��6q ~ q ~$5t 277t 113pw        sq ~#yZ��5q ~ q ~$5t 277t 125pw        sq ~#yZ��sq ~ q ~$5t 277t 127pw@$      sq ~#yZ�ڸq ~ q ~$5t 277t 133pw        sq ~#yZ��,q ~ q ~$5t 277t 30pw@$      sq ~#yZ��6q ~ q ~$5t 278t 103pw@$      sq ~#yZ��q ~ q ~$5t 278t 5pw@$      sq ~#yZ��q ~ q ~$5t 279t 61pw        sq ~#yZ��q ~ q ~$5t 279t 85pw@$      sq ~#yWŷ�q ~ q ~$5t 28t 26pw        sq ~#yW���q ~ q ~$5t 28t 66pw        sq ~#yW��eq ~ q ~$5t 28t 8pw@$      sq ~#yZ�)�q ~ q ~$5t 280t 103pw@$      sq ~#yZ�/lq ~ q ~$5t 280t 5pw@$      sq ~#yZ�3kq ~ q ~$5t 281t 7pw        sq ~#yZ�eq ~ q ~$5t 281t 85pw@$      sq ~#yZ���q ~ q ~$5t 282t 36pw        sq ~#yZ�	&q ~ q ~$5t 282t 85pw@$      sq ~#yZ��q ~ q ~$5t 283t 60pw        sq ~#yZ��q ~ q ~$5t 283t 85pw@$      sq ~#yZ�q ~ q ~$5t 283t 86pw@$      sq ~#yZ�8�q ~ q ~$5t 284t 103pw@$      sq ~#yZ�>pq ~ q ~$5t 284t 5pw@$      sq ~#yZ�	q ~ q ~$5t 285t 54pw@$      sq ~#yZ�K�q ~ q ~$5t 286t 137pw@$      sq ~#yZ�q ~ q ~$5t 286t 72pw@$      sq ~#yZ��q ~ q ~$5t 287t 54pw@5oz�G�sq ~#yZ��q ~ q ~$5t 288t 58pw        sq ~#yZ��q ~ q ~$5t 288t 85pw@$      sq ~#yZ�nq ~ q ~$5t 289t 73pw        sq ~#yZ�#mq ~ q ~$5t 289t 85pw@$      sq ~#yZ�#�q ~ q ~$5t 289t 86pw@$      sq ~#yWŻ�q ~ q ~$5t 29t 27pw@$      sq ~#yW��@q ~ q ~$5t 29t 75pw@$      sq ~#yZ�_q ~ q ~$5t 290t 21pw        sq ~#yZ��	q ~ q ~$5t 290t 7pw@$      sq ~#yZ���q ~ q ~$5t 291t 103pw@$      sq ~#yZ���q ~ q ~$5t 291t 5pw@$      sq ~#yZ�jcq ~ q ~$5t 292t 32pw@$      sq ~#yZ�r�q ~ q ~$5t 292t 58pw        sq ~#yZ�u�q ~ q ~$5t 293t 54pw@$      sq ~#yZ���q ~ q ~$5t 294t 112pw@$      sq ~#yZ��q ~ q ~$5t 294t 116pw        sq ~#yZ�n$q ~ q ~$5t 294t 22pw@$      sq ~#yZ��-q ~ q ~$5t 294t 90pw@$      sq ~#yZ��q ~ q ~$5t 295t 118pw        sq ~#yZ��,q ~ q ~$5t 295t 119pw@$      sq ~#yZ���q ~ q ~$5t 295t 120pw@$      sq ~#yZ���q ~ q ~$5t 295t 129pw        sq ~#yZ�ygq ~ q ~$5t 296t 32pw@$      sq ~#yZ��dq ~ q ~$5t 296t 68pw        sq ~#yZ��Kq ~ q ~$5t 297t 73pw        sq ~#yZ��Jq ~ q ~$5t 297t 85pw@$      sq ~#yZ��iq ~ q ~$5t 297t 86pw@$      sq ~#yZ��Pq ~ q ~$5t 298t 118pw@$      sq ~#yZ��q ~ q ~$5t 298t 120pw        sq ~#yZ��q ~ q ~$5t 298t 128pw        sq ~#yZ���q ~ q ~$5t 299t 121pw        sq ~#yZ���q ~ q ~$5t 299t 128pw@$      sq ~#yZ���q ~ q ~$5t 299t 96pw@$      sq ~#yW�.wq ~ q ~$5t 3t 3pw@$      sq ~#yW�/q ~ q ~$5t 3t 8pw@$      sq ~#yW��q ~ q ~$5t 30t 29pw        sq ~#yW�!3q ~ q ~$5t 30t 78pw@5oz�G�sq ~#yZ���q ~ q ~$5t 300t 137pw@$      sq ~#yZ�o'q ~ q ~$5t 300t 69pw@$      sq ~#yZ�rq ~ q ~$5t 300t 72pw        sq ~#yZ�f�q ~ q ~$5t 301t 32pw        sq ~#yZ�u�q ~ q ~$5t 301t 73pw@$      sq ~#yZ���q ~ q ~$5t 302t 103pw@$      sq ~#yZ��wq ~ q ~$5t 302t 5pw@$      sq ~#yZ��q ~ q ~$5t 303t 137pw@$      sq ~#yZ�}Rq ~ q ~$5t 303t 72pw@$      sq ~#yZ�~+q ~ q ~$5t 303t 79pw        sq ~#yZ�}q ~ q ~$5t 304t 60pw@$      sq ~#yZ��2q ~ q ~$5t 304t 73pw        sq ~#yZ���q ~ q ~$5t 305t 137pw@$      sq ~#yZ���q ~ q ~$5t 305t 72pw@$      sq ~#yZ��q ~ q ~$5t 306t 80pw@$      sq ~#yZ��q ~ q ~$5t 306t 92pw        sq ~#yZ�yrq ~ q ~$5t 307t 21pw        sq ~#yZ��tq ~ q ~$5t 307t 85pw@$      sq ~#yZ���q ~ q ~$5t 307t 86pw@$      sq ~#yZ��q ~ q ~$5t 308t 60pw        sq ~#yZ��5q ~ q ~$5t 308t 85pw@$      sq ~#yZ��Tq ~ q ~$5t 308t 86pw@$      sq ~#yZ���q ~ q ~$5t 309t 68pw        sq ~#yZ���q ~ q ~$5t 309t 73pw@$      sq ~#yW�Xq ~ q ~$5t 31t 125pw@$      sq ~#yW�[�q ~ q ~$5t 31t 133pw@$      sq ~#yW��q ~ q ~$5t 31t 30pw        sq ~#yZ�uq ~ q ~$5t 310t 103pw@$      sq ~#yZ�Tq ~ q ~$5t 310t 5pw@$      sq ~#yZ��q ~ q ~$5t 311t 122pw        sq ~#yZ��q ~ q ~$5t 311t 124pw@$      sq ~#yZ��q ~ q ~$5t 312t 54pw@F�U�i�sq ~#yZ�%:q ~ q ~$5t 313t 123pw        sq ~#yZ���q ~ q ~$5t 313t 84pw@$      sq ~#yZ��.q ~ q ~$5t 314t 54pw@$      sq ~#yZ�%:q ~ q ~$5t 315t 103pw@$      sq ~#yZ�+q ~ q ~$5t 315t 5pw@$      sq ~#yZ�0^q ~ q ~$5t 316t 122pw        sq ~#yZ�0�q ~ q ~$5t 316t 124pw@$      sq ~#yZ�4]q ~ q ~$5t 317t 124pw@$      sq ~#yZ�<<q ~ q ~$5t 318t 137pw@$      sq ~#yZ��q ~ q ~$5t 318t 69pw        sq ~#yZ�vq ~ q ~$5t 318t 72pw@$      sq ~#yZ�8q ~ q ~$5t 319t 60pw        sq ~#yZ�Uq ~ q ~$5t 319t 85pw@$      sq ~#yW��q ~ q ~$5t 32t 15pw        sq ~#yW�Y�q ~ q ~$5t 32t 3pw@$      sq ~#yW�Z>q ~ q ~$5t 32t 8pw@$      sq ~#yZ���q ~ q ~$5t 320t 103pw@$      sq ~#yZ���q ~ q ~$5t 320t 5pw@$      sq ~#yZ��q ~ q ~$5t 321t 111pw@$      sq ~#yZ�K�q ~ q ~$5t 321t 22pw@$      sq ~#yZ�fq ~ q ~$5t 321t 92pw        sq ~#yZ�f�q ~ q ~$5t 321t 97pw@$      sq ~#yZ�[q ~ q ~$5t 322t 54pw@$      sq ~#yZ��<q ~ q ~$5t 323t 120pw        sq ~#yZ��4q ~ q ~$5t 323t 128pw@5oz�G�sq ~#yZ�nq ~ q ~$5t 323t 96pw@5oz�G�sq ~#yZ�q4q ~ q ~$5t 324t 91pw@$      sq ~#yZ��q ~ q ~$5t 325t 130pw@5oz�G�sq ~#yZ�uqq ~ q ~$5t 325t 95pw@5oz�G�sq ~#yZ��q ~ q ~$5t 326t 137pw@$      sq ~#yZ�nkq ~ q ~$5t 326t 69pw@$      sq ~#yZ�r,q ~ q ~$5t 326t 79pw        sq ~#yZ��q ~ q ~$5t 327t 103pw@$      sq ~#yZ���q ~ q ~$5t 327t 5pw@$      sq ~#yZ���q ~ q ~$5t 328t 137pw@$      sq ~#yZ�u�q ~ q ~$5t 328t 69pw        sq ~#yZ�x�q ~ q ~$5t 328t 72pw@$      sq ~#yZ�y�q ~ q ~$5t 329t 68pw        sq ~#yZ���q ~ q ~$5t 329t 85pw@$      sq ~#yZ���q ~ q ~$5t 329t 86pw@$      sq ~#yW��q ~ q ~$5t 33t 27pw@$      sq ~#yW��q ~ q ~$5t 33t 33pw        sq ~#yW�,q ~ q ~$5t 33t 75pw@$      sq ~#yZ��(q ~ q ~$5t 330t 32pw        sq ~#yZ��Jq ~ q ~$5t 330t 85pw@$      sq ~#yZ��q ~ q ~$5t 331t 73pw        sq ~#yZ��q ~ q ~$5t 331t 85pw@$      sq ~#yZ�tq ~ q ~$5t 332t 137pw@5oz�G�sq ~#yZ���q ~ q ~$5t 332t 69pw@5oz�G�sq ~#yZ�Uq ~ q ~$5t 333t 126pw@@�鹙�sq ~#yZ��q ~ q ~$5t 334t 113pw        sq ~#yZ�q ~ q ~$5t 334t 114pw@$      sq ~#yZ�tq ~ q ~$5t 334t 117pw@$      sq ~#yZ�5q ~ q ~$5t 334t 127pw        sq ~#yZ��q ~ q ~$5t 335t 21pw@$      sq ~#yZ��q ~ q ~$5t 335t 61pw@$      sq ~#yZ�Sq ~ q ~$5t 335t 9pw        sq ~#yZ��q ~ q ~$5t 336t 103pw@$      sq ~#yZ��q ~ q ~$5t 336t 5pw@$      sq ~#yZ��lq ~ q ~$5t 337t 68pw        sq ~#yZ��q ~ q ~$5t 337t 85pw@5oz�G�sq ~#yZ��-q ~ q ~$5t 338t 68pw        sq ~#yZ��Rq ~ q ~$5t 338t 85pw@$      sq ~#yZ�(�q ~ q ~$5t 339t 137pw@$      sq ~#yZ���q ~ q ~$5t 339t 72pw@$      sq ~#yW�a%q ~ q ~$5t 34t 3pw@$      sq ~#yW� �q ~ q ~$5t 34t 34pw        sq ~#yW�a�q ~ q ~$5t 34t 8pw@$      sq ~#yZ�tq ~ q ~$5t 340t 119pw@$      sq ~#yZ�v�q ~ q ~$5t 340t 120pw@$      sq ~#yZ�v�q ~ q ~$5t 340t 121pw        sq ~#yZ�q ~ q ~$5t 341t 137pw@$      sq ~#yZ�GLq ~ q ~$5t 341t 72pw@$      sq ~#yZ�C�q ~ q ~$5t 342t 54pw@$      sq ~#yZ�V1q ~ q ~$5t 343t 91pw@$      sq ~#yZ�N�q ~ q ~$5t 344t 60pw        sq ~#yZ�V�q ~ q ~$5t 344t 85pw@@�鹙�sq ~#yZ���q ~ q ~$5t 345t 122pw        sq ~#yZ���q ~ q ~$5t 345t 124pw@i���sq ~#yZ�R�q ~ q ~$5t 345t 65pw@$      sq ~#yZ��q ~ q ~$5t 346t 103pw@$      sq ~#yZ���q ~ q ~$5t 346t 5pw@$      sq ~#yZ��q ~ q ~$5t 347t 105pw@$      sq ~#yZ�e�q ~ q ~$5t 348t 85pw@$      sq ~#yZ�e�q ~ q ~$5t 348t 86pw@$      sq ~#yZ��q ~ q ~$5t 349t 137pw@$      sq ~#yZ�blq ~ q ~$5t 349t 69pw        sq ~#yZ�eTq ~ q ~$5t 349t 72pw@$      sq ~#yW�$�q ~ q ~$5t 35t 35pw        sq ~#yW�e�q ~ q ~$5t 35t 8pw@$      sq ~#yZ��Mq ~ q ~$5t 350t 91pw@-����ŀsq ~#yZ��gq ~ q ~$5t 351t 54pw@$      sq ~#yZ��(q ~ q ~$5t 352t 54pw@$      sq ~#yZ���q ~ q ~$5t 353t 137pw@$      sq ~#yZ��-q ~ q ~$5t 353t 72pw@$      sq ~#yZ��q ~ q ~$5t 353t 79pw        sq ~#yZ���q ~ q ~$5t 354t 103pw@$      sq ~#yZ���q ~ q ~$5t 354t 5pw@$      sq ~#yZ��gq ~ q ~$5t 355t 14pw        sq ~#yZ���q ~ q ~$5t 355t 85pw@$      sq ~#yZ�Ҏq ~ q ~$5t 356t 85pw@$      sq ~#yZ�ҭq ~ q ~$5t 356t 86pw@$      sq ~#yZ� �q ~ q ~$5t 356t 9pw        sq ~#yZ�	�q ~ q ~$5t 357t 137pw@$      sq ~#yZ��1q ~ q ~$5t 357t 72pw@$      sq ~#yZ��q ~ q ~$5t 358t 103pw@$      sq ~#yZ��q ~ q ~$5t 358t 5pw@$      sq ~#yZ�yq ~ q ~$5t 359t 137pw@5oz�G�sq ~#yZ�ٳq ~ q ~$5t 359t 72pw@5oz�G�sq ~#yW�$�q ~ q ~$5t 36t 26pw@5oz�G�sq ~#yW�(q ~ q ~$5t 36t 33pw        sq ~#yZ�_�q ~ q ~$5t 360t 122pw@$      sq ~#yZ�_�q ~ q ~$5t 360t 124pw@$      sq ~#yZ�(�q ~ q ~$5t 360t 65pw        sq ~#yZ�\q ~ q ~$5t 361t 103pw@$      sq ~#yZ�a�q ~ q ~$5t 361t 5pw@$      sq ~#yZ�j�q ~ q ~$5t 362t 132pw@5oz�G�sq ~#yZ�oRq ~ q ~$5t 363t 137pw@$      sq ~#yZ�4�q ~ q ~$5t 363t 69pw        sq ~#yZ�7�q ~ q ~$5t 363t 72pw@$      sq ~#yZ�4	q ~ q ~$5t 364t 54pw@ �̾�,sq ~#yZ�kq ~ q ~$5t 365t 103pw@@�鹙�sq ~#yZ�p�q ~ q ~$5t 365t 5pw@@�鹙�sq ~#yZ�;�q ~ q ~$5t 366t 54pw@$      sq ~#yZ�r�q ~ q ~$5t 367t 105pw@$      sq ~#yZ��>q ~ q ~$5t 368t 130pw@$      sq ~#yZ�R0q ~ q ~$5t 368t 95pw@$      sq ~#yZ���q ~ q ~$5t 369t 137pw@%��9�}qsq ~#yZ�Nq ~ q ~$5t 369t 72pw@$      sq ~#yW�lq ~ q ~$5t 37t 0pw        sq ~#yW�lhq ~ q ~$5t 37t 3pw@#��吢sq ~#yW�mq ~ q ~$5t 37t 8pw@$      sq ~#yZ��dq ~ q ~$5t 370t 54pw@$      sq ~#yZ��pq ~ q ~$5t 371t 103pw@$      sq ~#yZ��Oq ~ q ~$5t 371t 5pw@$      sq ~#yZ���q ~ q ~$5t 372t 124pw@$      sq ~#yZ���q ~ q ~$5t 373t 54pw@&'��5V�sq ~#yZ��rq ~ q ~$5t 374t 137pw@$      sq ~#yZ���q ~ q ~$5t 374t 69pw        sq ~#yZ���q ~ q ~$5t 374t 72pw@$      sq ~#yZ��)q ~ q ~$5t 375t 54pw@$      sq ~#yZ��5q ~ q ~$5t 376t 103pw@$      sq ~#yZ��q ~ q ~$5t 376t 5pw@$      sq ~#yZ���q ~ q ~$5t 377t 54pw@$      sq ~#yZ��q ~ q ~$5t 378t 103pw@$      sq ~#yZ��q ~ q ~$5t 378t 5pw@$      sq ~#yZ��7q ~ q ~$5t 379t 137pw@$      sq ~#yZ���q ~ q ~$5t 379t 69pw        sq ~#yZ��qq ~ q ~$5t 379t 72pw@$      sq ~#yW�j+q ~ q ~$5t 38t 100pw@$      sq ~#yW�0q ~ q ~$5t 38t 37pw        sq ~#yW�?;q ~ q ~$5t 38t 78pw        sq ~#yW�B�q ~ q ~$5t 38t 87pw@$      sq ~#yW�F"q ~ q ~$5t 38t 93pw@$      sq ~#yZ��q ~ q ~$5t 380t 54pw@$      sq ~#yZ�D�q ~ q ~$5t 381t 103pw@$      sq ~#yZ�J�q ~ q ~$5t 381t 5pw@$      sq ~#yZ�H�q ~ q ~$5t 382t 103pw@$      sq ~#yZ�Noq ~ q ~$5t 382t 5pw@$      sq ~#yZ�q ~ q ~$5t 383t 54pw@$      sq ~#yZ��q ~ q ~$5t 384t 54pw@$      sq ~#yZ�S�q ~ q ~$5t 385t 103pw@5oz�G�sq ~#yZ�Y�q ~ q ~$5t 385t 5pw@5oz�G�sq ~#yZ�$Iq ~ q ~$5t 386t 54pw@5oz�G�sq ~#yZ�f;q ~ q ~$5t 387t 130pw@$      sq ~#yZ�7-q ~ q ~$5t 387t 95pw@$      sq ~#yZ�_q ~ q ~$5t 388t 103pw@$      sq ~#yZ�d�q ~ q ~$5t 388t 5pw@$      sq ~#yZ�jxq ~ q ~$5t 389t 124pw@$      sq ~#yW�3�q ~ q ~$5t 39t 38pw        sq ~#yW�t�q ~ q ~$5t 39t 8pw@$      sq ~#yZ���q ~ q ~$5t 390t 91pw@$      sq ~#yZ��.q ~ q ~$5t 391t 103pw@5oz�G�sq ~#yZ��q ~ q ~$5t 391t 5pw@5oz�G�sq ~#yZ���q ~ q ~$5t 392t 103pw@$      sq ~#yZ���q ~ q ~$5t 392t 5pw@$      sq ~#yZ���q ~ q ~$5t 393t 103pw@5oz�G�sq ~#yZ�Əq ~ q ~$5t 393t 5pw@5oz�G�sq ~#yZ��qq ~ q ~$5t 394t 103pw@$      sq ~#yZ��Pq ~ q ~$5t 394t 5pw@$      sq ~#yZ��2q ~ q ~$5t 395t 103pw@$      sq ~#yZ��q ~ q ~$5t 395t 5pw@$      sq ~#yZ�ײq ~ q ~$5t 396t 137pw@F�U�i�sq ~#yZ��q ~ q ~$5t 396t 69pw@F�U�i�sq ~#yZ���q ~ q ~$5t 396t 72pw        sq ~#yZ��iq ~ q ~$5t 397t 54pw@5oz�G�sq ~#yZ��4q ~ q ~$5t 398t 137pw@$      sq ~#yZ���q ~ q ~$5t 398t 69pw@$      sq ~#yZ���q ~ q ~$5t 399t 137pw@$      sq ~#yZ��/q ~ q ~$5t 399t 72pw@$      sq ~#yZ��q ~ q ~$5t 399t 79pw        sq ~#yW�28q ~ q ~$5t 4t 3pw@&��}�sq ~#yW�2Wq ~ q ~$5t 4t 4pw        sq ~#yW��Mq ~ q ~$5t 4t 42pw���]=���sq ~#yW�2�q ~ q ~$5t 4t 8pw@$      sq ~#yWƆ�q ~ q ~$5t 40t 39pw        sq ~#yW��q ~ q ~$5t 40t 8pw@5v��n�sq ~#yZ��Lq ~ q ~$5t 400t 54pw@$      sq ~#yZ��Xq ~ q ~$5t 401t 103pw@$      sq ~#yZ��7q ~ q ~$5t 401t 5pw@$      sq ~#yZ���q ~ q ~$5t 402t 137pw@$      sq ~#yZ��q ~ q ~$5t 402t 72pw@$      sq ~#yZ��<q ~ q ~$5t 403t 134pw@5oz�G�sq ~#yZ�Ͽq ~ q ~$5t 404t 132pw@$      sq ~#yZ��q ~ q ~$5t 405t 54pw@$      sq ~#yZ��Aq ~ q ~$5t 406t 132pw@$      sq ~#yZ��q ~ q ~$5t 407t 132pw@$      sq ~#yZ��^q ~ q ~$5t 408t 137pw@$      sq ~#yZ���q ~ q ~$5t 408t 72pw@$      sq ~#yZ��`q ~ q ~$5t 409t 103pw@$      sq ~#yZ��?q ~ q ~$5t 409t 5pw@$      sq ~#yWƂ2q ~ q ~$5t 41t 13pw        sq ~#yWƉ�q ~ q ~$5t 41t 34pw@$      sq ~#yWƍuq ~ q ~$5t 41t 43pw        sq ~#yZ�5q ~ q ~$5t 410t 132pw@$      sq ~#yZ�-�q ~ q ~$5t 411t 103pw@5oz�G�sq ~#yZ�3�q ~ q ~$5t 411t 5pw@5oz�G�sq ~#yZ�1�q ~ q ~$5t 412t 105pw@$      sq ~#yZ��q ~ q ~$5t 413t 54pw@$      sq ~#yZ��q ~ q ~$5t 414t 54pw@$      sq ~#yZ�<�q ~ q ~$5t 415t 103pw@5oz�G�sq ~#yZ�B�q ~ q ~$5t 415t 5pw@5oz�G�sq ~#yZ�1q ~ q ~$5t 416t 54pw@$      sq ~#yZ��q ~ q ~$5t 417t 54pw@$      sq ~#yZ��q ~ q ~$5t 418t 54pw@$      sq ~#yZ�V�q ~ q ~$5t 419t 130pw@$      sq ~#yZ�'�q ~ q ~$5t 419t 95pw@$      sq ~#yW��q ~ q ~$5t 42t 3pw@5oz�G�sq ~#yWƐ�q ~ q ~$5t 42t 40pw        sq ~#yW�Νq ~ q ~$5t 42t 8pw@5oz�G�sq ~#yZ�k
q ~ q ~$5t 420t 54pw@@�鹙�sq ~#yZ��Tq ~ q ~$5t 421t 105pw@5oz�G�sq ~#yZ�r�q ~ q ~$5t 422t 54pw@$      sq ~#yZ�vMq ~ q ~$5t 423t 54pw@5oz�G�sq ~#yZ�zq ~ q ~$5t 424t 54pw@$      sq ~#yZ���q ~ q ~$5t 425t 135pw@@�鹙�sq ~#yZ���q ~ q ~$5t 426t 54pw@$      sq ~#yZ��<q ~ q ~$5t 427t 136pw@@�鹙�sq ~#yZ��q ~ q ~$5t 428t 54pw@5oz�G�sq ~#yZ��+q ~ q ~$5t 429t 29pw        sq ~#yZ���q ~ q ~$5t 429t 93pw@�iu��sq ~#yWƍ�q ~ q ~$5t 43t 27pw@$�g\oQsq ~#yWƔ�q ~ q ~$5t 43t 41pw        sq ~#yWƕ5q ~ q ~$5t 43t 45pw        sq ~#yWƠxq ~ q ~$5t 43t 75pw@$      sq ~#yZ�ԃq ~ q ~$5t 430t 27pw?��C1S_sq ~#yZ�tq ~ q ~$5t 430t 4pw        sq ~#yZ��jq ~ q ~$5t 430t 42pw@j ���sq ~#yZ��Cq ~ q ~$5t 430t 49pw@8�q;Hsq ~#yZ��q ~ q ~$5t 430t 8pw?��$*pRsq ~#yZ�q ~ q ~$5t 431t 124pw?��2Q�v�sq ~#yZ��
q ~ q ~$5t 431t 65pw        sq ~#yZ�!�q ~ q ~$5t 432t 124pw@�xJdGsq ~#yZ���q ~ q ~$5t 433t 20pw        sq ~#yZ��q ~ q ~$5t 433t 42pw@$��D��asq ~#yZ��Lq ~ q ~$5t 434t 77pw        sq ~#yZ�'�q ~ q ~$5t 434t 8pw@�<�/ssq ~#yZ���q ~ q ~$5t 435t 74pw        sq ~#yZ��q ~ q ~$5t 435t 99pw?��s��֓sq ~#yZ�oq ~ q ~$5t 436t 98pw        sq ~#yZ��q ~ q ~$5t 436t 99pw?��s��֓sq ~#yZ���q ~ q ~$5t 437t 39pw        sq ~#yZ���q ~ q ~$5t 437t 42pw@sw�:sq ~#yZ�8]q ~ q ~$5t 438t 124pw@���Nsq ~#yZ�Qq ~ q ~$5t 438t 65pw        sq ~#yWƐ�q ~ q ~$5t 44t 21pw        sq ~#yWƧ�q ~ q ~$5t 44t 85pw@5oz�G�sq ~#yW��&q ~ q ~$5t 45t 2pw@5oz�G�sq ~#yWƔ�q ~ q ~$5t 45t 20pw@5oz�G�sq ~#yWƜZq ~ q ~$5t 45t 42pw        sq ~#yWƠq ~ q ~$5t 46t 42pw@$      sq ~#yWƠYq ~ q ~$5t 46t 44pw        sq ~#yWƘ�q ~ q ~$5t 47t 13pw        sq ~#yWƮ�q ~ q ~$5t 47t 70pw@$      sq ~#yW��q ~ q ~$5t 48t 3pw@$�g\oIsq ~#yWƤq ~ q ~$5t 48t 34pw        sq ~#yW��#q ~ q ~$5t 48t 8pw@$      sq ~#yWƠ�q ~ q ~$5t 49t 17pw@$      sq ~#yWƫ�q ~ q ~$5t 49t 46pw        sq ~#yW�0Xq ~ q ~$5t 5t 103pw@5oz�G�sq ~#yW�67q ~ q ~$5t 5t 5pw@5oz�G�sq ~#yW��kq ~ q ~$5t 50t 18pw        sq ~#yW�;zq ~ q ~$5t 50t 8pw@$      sq ~#yW���q ~ q ~$5t 51t 20pw        sq ~#yW�?;q ~ q ~$5t 51t 8pw@$      sq ~#yW�0q ~ q ~$5t 52t 48pw        sq ~#yW�B�q ~ q ~$5t 52t 8pw@$      sq ~#yW�F"q ~ q ~$5t 53t 3pw@5oz�G�sq ~#yW�
q ~ q ~$5t 53t 49pw        sq ~#yW�q ~ q ~$5t 53t 53pw        sq ~#yW�F�q ~ q ~$5t 53t 8pw@5oz�G�sq ~#yW��q ~ q ~$5t 54t 12pw        sq ~#yW�J~q ~ q ~$5t 54t 8pw@$      sq ~#yW�0q ~ q ~$5t 55t 18pw        sq ~#yW�N?q ~ q ~$5t 55t 8pw@$      sq ~#yW�Q�q ~ q ~$5t 56t 4pw@5oz�G�sq ~#yW��q ~ q ~$5t 56t 50pw        sq ~#yW� q ~ q ~$5t 56t 75pw        sq ~#yW� Xq ~ q ~$5t 56t 77pw        sq ~#yW�O(q ~ q ~$5t 57t 100pw        sq ~#yW�OGq ~ q ~$5t 57t 101pw@$      sq ~#yW�Pq ~ q ~$5t 57t 107pw@$      sq ~#yW��q ~ q ~$5t 57t 29pw@$      sq ~#yW��q ~ q ~$5t 57t 51pw        sq ~#yW�'?q ~ q ~$5t 57t 82pw@$      sq ~#yW�+�q ~ q ~$5t 57t 99pw        sq ~#yW�Yq ~ q ~$5t 58t 45pw@$      sq ~#yW��q ~ q ~$5t 58t 52pw        sq ~#yW��q ~ q ~$5t 59t 26pw        sq ~#yW��q ~ q ~$5t 59t 27pw��N>)L�&sq ~#yW��q ~ q ~$5t 59t 42pw@�e��'�sq ~#yW���q ~ q ~$5t 6t 15pw        sq ~#yW���q ~ q ~$5t 6t 27pw@$      sq ~#yW�:q ~ q ~$5t 6t 6pw        sq ~#yW�oq ~ q ~$5t 6t 75pw@$      sq ~#yWƮ�q ~ q ~$5t 60t 0pw        sq ~#yW�gmq ~ q ~$5t 60t 15pw@$      sq ~#yW�klq ~ q ~$5t 60t 27pw��N>)L�&sq ~#yW�rSq ~ q ~$5t 60t 42pw@�e��'�sq ~#yW�zq ~ q ~$5t 61t 54pw@$      sq ~#yW�}�q ~ q ~$5t 62t 55pw        sq ~#yW�~oq ~ q ~$5t 62t 59pw@5oz�G�sq ~#yW�v�q ~ q ~$5t 63t 27pw@$      sq ~#yWǁ�q ~ q ~$5t 63t 56pw        sq ~#yWǉ6q ~ q ~$5t 63t 75pw@$      sq ~#yW�v�q ~ q ~$5t 64t 19pw        sq ~#yWƾBq ~ q ~$5t 64t 3pw@$      sq ~#yWƾ�q ~ q ~$5t 64t 8pw@$      sq ~#yW�~1q ~ q ~$5t 65t 27pw@$      sq ~#yWǉtq ~ q ~$5t 65t 57pw        sq ~#yWǐ�q ~ q ~$5t 65t 75pw@$      sq ~#yW�}�q ~ q ~$5t 66t 12pw        sq ~#yW���q ~ q ~$5t 66t 3pw@$      sq ~#yW��_q ~ q ~$5t 66t 8pw@$      sq ~#yWǁ�q ~ q ~$5t 67t 14pw@$      sq ~#yWǄ�q ~ q ~$5t 67t 21pw@$      sq ~#yWǑq ~ q ~$5t 67t 58pw        sq ~#yW��Fq ~ q ~$5t 68t 3pw@5oz�G�sq ~#yWǔ;q ~ q ~$5t 68t 53pw        sq ~#yW���q ~ q ~$5t 68t 8pw@5oz�G�sq ~#yWǘ�q ~ q ~$5t 69t 58pw������c�sq ~#yWǣ}q ~ q ~$5t 69t 85pw@$      sq ~#yW��q ~ q ~$5t 7t 60pw@$      sq ~#yW�=�q ~ q ~$5t 7t 7pw        sq ~#yW���q ~ q ~$5t 70t 60pw        sq ~#yW��q ~ q ~$5t 70t 73pw@$      sq ~#yW��q ~ q ~$5t 71t 11pw        sq ~#yW��Wq ~ q ~$5t 71t 93pw@5oz�G�sq ~#yW�+q ~ q ~$5t 72t 3pw@5oz�G�sq ~#yW��q ~ q ~$5t 72t 41pw        sq ~#yW�+�q ~ q ~$5t 72t 8pw@5oz�G�sq ~#yW��q ~ q ~$5t 73t 15pw        sq ~#yW��-q ~ q ~$5t 73t 28pw@$      sq ~#yW�2�q ~ q ~$5t 74t 3pw@@�鹙�sq ~#yW��xq ~ q ~$5t 74t 40pw        sq ~#yW�3<q ~ q ~$5t 74t 8pw@@�鹙�sq ~#yW��9q ~ q ~$5t 75t 40pw        sq ~#yW�6�q ~ q ~$5t 75t 8pw@$      sq ~#yW�7q ~ q ~$5t 76t 54pw@$      sq ~#yW�=�q ~ q ~$5t 77t 1pw@$      sq ~#yW�6q ~ q ~$5t 77t 56pw@$      sq ~#yW�>q ~ q ~$5t 77t 8pw        sq ~#yW��q ~ q ~$5t 78t 21pw        sq ~#yW�q ~ q ~$5t 78t 85pw@$      sq ~#yW�:q ~ q ~$5t 78t 86pw@$      sq ~#yW���q ~ q ~$5t 79t 16pw        sq ~#yW��q ~ q ~$5t 79t 27pw@$      sq ~#yW�q ~ q ~$5t 79t 75pw@$      sq ~#yW�@�q ~ q ~$5t 8t 0pw@@�鹙�sq ~#yW�A�q ~ q ~$5t 8t 8pw        sq ~#yW�W�q ~ q ~$5t 80t 36pw        sq ~#yW�jrq ~ q ~$5t 80t 85pw@$      sq ~#yW�S�q ~ q ~$5t 81t 13pw        sq ~#yW�W�q ~ q ~$5t 81t 25pw@$      sq ~#yWǟ~q ~ q ~$5t 82t 3pw@$      sq ~#yW�_�q ~ q ~$5t 82t 39pw        sq ~#yWǠq ~ q ~$5t 82t 8pw@$      sq ~#yW�[nq ~ q ~$5t 83t 15pw        sq ~#yW�i�q ~ q ~$5t 83t 50pw@$      sq ~#yWǧ q ~ q ~$5t 84t 3pw@@�鹙�sq ~#yW�n3q ~ q ~$5t 84t 55pw        sq ~#yWǧ�q ~ q ~$5t 84t 8pw@@�鹙�sq ~#yWǪ�q ~ q ~$5t 85t 3pw@$      sq ~#yW�m�q ~ q ~$5t 85t 40pw        sq ~#yWǫ\q ~ q ~$5t 85t 8pw@$      sq ~#yW�j�q ~ q ~$5t 86t 26pw@5oz�G�sq ~#yW�u�q ~ q ~$5t 86t 57pw        sq ~#yW�|�q ~ q ~$5t 87t 61pw        sq ~#yWȀ�q ~ q ~$5t 87t 73pw@$      sq ~#yW�q�q ~ q ~$5t 88t 23pw        sq ~#yW�r2q ~ q ~$5t 88t 27pw@$      sq ~#yWȄ�q ~ q ~$5t 88t 75pw@$      sq ~#yWǹ�q ~ q ~$5t 89t 3pw@$      sq ~#yW�y�q ~ q ~$5t 89t 38pw        sq ~#yWǺ`q ~ q ~$5t 89t 8pw@$      sq ~#yW�sq ~ q ~$5t 9t 85pw@$      sq ~#yW��q ~ q ~$5t 9t 86pw@$      sq ~#yW�E�q ~ q ~$5t 9t 9pw        sq ~#yW�Ϗq ~ q ~$5t 90t 43pw@$      sq ~#yW�Ϯq ~ q ~$5t 90t 44pw        sq ~#yW�
�q ~ q ~$5t 91t 104pw@$      sq ~#yW���q ~ q ~$5t 91t 51pw@$      sq ~#yW�ڳq ~ q ~$5t 91t 62pw        sq ~#yW��q ~ q ~$5t 91t 93pw        sq ~#yW�Ϗq ~ q ~$5t 92t 23pw@5oz�G�sq ~#yW��q ~ q ~$5t 92t 55pw        sq ~#yW��0q ~ q ~$5t 93t 34pw        sq ~#yW�ޓq ~ q ~$5t 93t 53pw@$      sq ~#yW��
q ~ q ~$5t 94t 19pw@$      sq ~#yW��0q ~ q ~$5t 94t 24pw        sq ~#yW��5q ~ q ~$5t 94t 52pw@$      sq ~#yW���q ~ q ~$5t 95t 63pw        sq ~#yW��q ~ q ~$5t 95t 8pw@$      sq ~#yW��5q ~ q ~$5t 96t 32pw@$      sq ~#yW��:q ~ q ~$5t 96t 60pw        sq ~#yW�$�q ~ q ~$5t 97t 112pw@$      sq ~#yW��wq ~ q ~$5t 97t 64pw        sq ~#yW��>q ~ q ~$5t 97t 90pw@$      sq ~#yW�,cq ~ q ~$5t 98t 124pw@i���sq ~#yW��Wq ~ q ~$5t 98t 65pw        sq ~#yW���q ~ q ~$5t 99t 61pw        sq ~#yW� �q ~ q ~$5t 99t 85pw@$      sq ~#yW� �q ~ q ~$5t 99t 86pw@$      q ~#~w?�      sq ~#ye��q ~ t TMPt 0ppw?�ELE.tsq ~#ye���q ~ q ~00t 1ppw        sq ~#ye�A>q ~ q ~00t 10ppw        sq ~#yh�L�q ~ q ~00t 100ppw        sq ~#yh�PQq ~ q ~00t 101ppw        sq ~#yh�Tq ~ q ~00t 102ppw        sq ~#yh�W�q ~ q ~00t 103ppw        sq ~#yh�[�q ~ q ~00t 104ppw        sq ~#yh�_Uq ~ q ~00t 105ppw        sq ~#yh�cq ~ q ~00t 106ppw        sq ~#yh�f�q ~ q ~00t 107ppw?��b���Tsq ~#yh�j�q ~ q ~00t 108ppw        sq ~#yh�nYq ~ q ~00t 109ppw        sq ~#ye�D�q ~ q ~00t 11ppw        sq ~#yh���q ~ q ~00t 110ppw        sq ~#yh�İq ~ q ~00t 111ppw        sq ~#yh��qq ~ q ~00t 112ppw        sq ~#yh��2q ~ q ~00t 113ppw        sq ~#yh���q ~ q ~00t 114ppw        sq ~#yh�Ӵq ~ q ~00t 115ppw        sq ~#yh��uq ~ q ~00t 116ppw        sq ~#yh��6q ~ q ~00t 117ppw        sq ~#yh���q ~ q ~00t 118ppw        sq ~#yh��q ~ q ~00t 119ppw        sq ~#ye�H�q ~ q ~00t 12ppw        sq ~#yh�5Nq ~ q ~00t 120ppw        sq ~#yh�9q ~ q ~00t 121ppw        sq ~#yh�<�q ~ q ~00t 122ppw        sq ~#yh�@�q ~ q ~00t 123ppw        sq ~#yh�DRq ~ q ~00t 124ppw?��h%�-sq ~#yh�Hq ~ q ~00t 125ppw        sq ~#yh�K�q ~ q ~00t 126ppw        sq ~#yh�O�q ~ q ~00t 127ppw        sq ~#yh�SVq ~ q ~00t 128ppw        sq ~#yh�Wq ~ q ~00t 129ppw        sq ~#ye�L�q ~ q ~00t 13ppw        sq ~#yh���q ~ q ~00t 130ppw        sq ~#yh��nq ~ q ~00t 131ppw        sq ~#yh��/q ~ q ~00t 132ppw        sq ~#yh���q ~ q ~00t 133ppw        sq ~#yh���q ~ q ~00t 134ppw        sq ~#yh��rq ~ q ~00t 135ppw        sq ~#yh��3q ~ q ~00t 136ppw        sq ~#yh���q ~ q ~00t 137ppw?�Z�o���sq ~#ye�PBq ~ q ~00t 14ppw        sq ~#ye�Tq ~ q ~00t 15ppw        sq ~#ye�W�q ~ q ~00t 16ppw        sq ~#ye�[�q ~ q ~00t 17ppw        sq ~#ye�_Fq ~ q ~00t 18ppw        sq ~#ye�cq ~ q ~00t 19ppw        sq ~#ye��q ~ q ~00t 2ppw        sq ~#yeص�q ~ q ~00t 20ppw        sq ~#yeع^q ~ q ~00t 21ppw        sq ~#yeؽq ~ q ~00t 22ppw        sq ~#ye���q ~ q ~00t 23ppw        sq ~#ye�ġq ~ q ~00t 24ppw        sq ~#ye��bq ~ q ~00t 25ppw        sq ~#ye��#q ~ q ~00t 26ppw?���Mo�sq ~#ye���q ~ q ~00t 27ppw���3�sq ~#ye�ӥq ~ q ~00t 28ppw        sq ~#ye��fq ~ q ~00t 29ppw        sq ~#ye�Rq ~ q ~00t 3ppw���T����sq ~#ye�)�q ~ q ~00t 30ppw        sq ~#ye�-�q ~ q ~00t 31ppw        sq ~#ye�1~q ~ q ~00t 32ppw        sq ~#ye�5?q ~ q ~00t 33ppw        sq ~#ye�9 q ~ q ~00t 34ppw        sq ~#ye�<�q ~ q ~00t 35ppw        sq ~#ye�@�q ~ q ~00t 36ppw        sq ~#ye�DCq ~ q ~00t 37ppw        sq ~#ye�Hq ~ q ~00t 38ppw        sq ~#ye�K�q ~ q ~00t 39ppw        sq ~#ye�
q ~ q ~00t 4ppw        sq ~#yeٞ[q ~ q ~00t 40ppw        sq ~#ye٢q ~ q ~00t 41ppw        sq ~#ye٥�q ~ q ~00t 42ppw?���X�Fsq ~#ye٩�q ~ q ~00t 43ppw        sq ~#ye٭_q ~ q ~00t 44ppw        sq ~#yeٱ q ~ q ~00t 45ppw        sq ~#yeٴ�q ~ q ~00t 46ppw        sq ~#yeٸ�q ~ q ~00t 47ppw        sq ~#yeټcq ~ q ~00t 48ppw        sq ~#ye��$q ~ q ~00t 49ppw��>h3��sq ~#ye��q ~ q ~00t 5ppw        sq ~#ye��q ~ q ~00t 50ppw        sq ~#ye�{q ~ q ~00t 51ppw        sq ~#ye�<q ~ q ~00t 52ppw        sq ~#ye��q ~ q ~00t 53ppw        sq ~#ye�!�q ~ q ~00t 54ppw?�\����usq ~#ye�%q ~ q ~00t 55ppw        sq ~#ye�)@q ~ q ~00t 56ppw        sq ~#ye�-q ~ q ~00t 57ppw        sq ~#ye�0�q ~ q ~00t 58ppw�������sq ~#ye�4�q ~ q ~00t 59ppw        sq ~#ye��q ~ q ~00t 6ppw        sq ~#yeڇq ~ q ~00t 60ppw        sq ~#yeڊ�q ~ q ~00t 61ppw        sq ~#yeڎ�q ~ q ~00t 62ppw        sq ~#yeڒ\q ~ q ~00t 63ppw        sq ~#yeږq ~ q ~00t 64ppw��z©8sq ~#yeڙ�q ~ q ~00t 65ppw        sq ~#yeڝ�q ~ q ~00t 66ppw��Ŋ��sq ~#yeڡ`q ~ q ~00t 67ppw        sq ~#yeڥ!q ~ q ~00t 68ppw        sq ~#yeڨ�q ~ q ~00t 69ppw?��E��|`sq ~#ye�Vq ~ q ~00t 7ppw        sq ~#ye��xq ~ q ~00t 70ppw        sq ~#ye��9q ~ q ~00t 71ppw�΀�%R��sq ~#ye��q ~ q ~00t 72ppw?�a*0psq ~#ye��q ~ q ~00t 73ppw        sq ~#ye�
|q ~ q ~00t 74ppw        sq ~#ye�=q ~ q ~00t 75ppw        sq ~#ye��q ~ q ~00t 76ppw        sq ~#ye��q ~ q ~00t 77ppw        sq ~#ye��q ~ q ~00t 78ppw        sq ~#ye�Aq ~ q ~00t 79ppw        sq ~#ye�q ~ q ~00t 8ppw?ْR���sq ~#ye�o�q ~ q ~00t 80ppw        sq ~#ye�s�q ~ q ~00t 81ppw        sq ~#ye�wYq ~ q ~00t 82ppw        sq ~#ye�{q ~ q ~00t 83ppw        sq ~#ye�~�q ~ q ~00t 84ppw        sq ~#yeۂ�q ~ q ~00t 85ppw?�g�-�usq ~#yeۆ]q ~ q ~00t 86ppw        sq ~#yeۊq ~ q ~00t 87ppw        sq ~#yeۍ�q ~ q ~00t 88ppw        sq ~#yeۑ�q ~ q ~00t 89ppw��z©8sq ~#ye��q ~ q ~00t 9ppw        sq ~#ye��6q ~ q ~00t 90ppw        sq ~#ye���q ~ q ~00t 91ppw?��b���Gsq ~#ye��q ~ q ~00t 92ppw�΀�%R��sq ~#ye��yq ~ q ~00t 93ppw?��)��sq ~#ye��:q ~ q ~00t 94ppw        sq ~#ye���q ~ q ~00t 95ppw        sq ~#ye���q ~ q ~00t 96ppw        sq ~#ye��}q ~ q ~00t 97ppw�΀�%R��sq ~#ye�>q ~ q ~00t 98ppw        sq ~#ye��q ~ q ~00t 99ppw?���9+��q ~#zw?�      sq ~#y{H�q ~ t XEMEt 0ppw@$      sq ~#y{H��q ~ q ~1Et 1ppw@$      sq ~#y{^�0q ~ q ~1Et 10ppw@$      sq ~#y~��q ~ q ~1Et 100ppw@$      sq ~#y~�Cq ~ q ~1Et 101ppw@'���@nsq ~#y~q ~ q ~1Et 102ppw@;�뤍sq ~#y~�q ~ q ~1Et 103ppw@$      sq ~#y~�q ~ q ~1Et 104ppw@$      sq ~#y~Gq ~ q ~1Et 105ppw@%��9�}isq ~#y~q ~ q ~1Et 106ppw@$      sq ~#y~�q ~ q ~1Et 107ppw@$      sq ~#y~�q ~ q ~1Et 108ppw@$      sq ~#y~Kq ~ q ~1Et 109ppw@$      sq ~#y{^��q ~ q ~1Et 11ppw@$      sq ~#y~m�q ~ q ~1Et 110ppw@$      sq ~#y~q�q ~ q ~1Et 111ppw@$      sq ~#y~ucq ~ q ~1Et 112ppw@#��吢sq ~#y~y$q ~ q ~1Et 113ppw@)r�|��sq ~#y~|�q ~ q ~1Et 114ppw@$      sq ~#y~��q ~ q ~1Et 115ppw@$      sq ~#y~�gq ~ q ~1Et 116ppw@$      sq ~#y~�(q ~ q ~1Et 117ppw@$      sq ~#y~��q ~ q ~1Et 118ppw@$      sq ~#y~��q ~ q ~1Et 119ppw@$      sq ~#y{^��q ~ q ~1Et 12ppw@$      sq ~#y~�@q ~ q ~1Et 120ppw@$      sq ~#y~�q ~ q ~1Et 121ppw@'���@nsq ~#y~��q ~ q ~1Et 122ppw@$      sq ~#y~�q ~ q ~1Et 123ppw@"
\�Hq�sq ~#y~�Dq ~ q ~1Et 124ppw@$      sq ~#y~�q ~ q ~1Et 125ppw@$      sq ~#y~��q ~ q ~1Et 126ppw@%U�i�g�sq ~#y~��q ~ q ~1Et 127ppw@$      sq ~#y~ Hq ~ q ~1Et 128ppw@$      sq ~#y~	q ~ q ~1Et 129ppw@$      sq ~#y{^�sq ~ q ~1Et 13ppw@$      sq ~#y~V�q ~ q ~1Et 130ppw@$      sq ~#y~Z`q ~ q ~1Et 131ppw@$      sq ~#y~^!q ~ q ~1Et 132ppw@$      sq ~#y~a�q ~ q ~1Et 133ppw@$      sq ~#y~e�q ~ q ~1Et 134ppw@$      sq ~#y~idq ~ q ~1Et 135ppw@#]<6(��sq ~#y~m%q ~ q ~1Et 136ppw@$      sq ~#y~p�q ~ q ~1Et 137ppw@$      sq ~#y~t�q ~ q ~1Et 138ppw@$      sq ~#y~xhq ~ q ~1Et 139ppw@$      sq ~#y{^�4q ~ q ~1Et 14ppw@$      sq ~#y~��q ~ q ~1Et 140ppw@$      sq ~#y~οq ~ q ~1Et 141ppw@$      sq ~#y~Ҁq ~ q ~1Et 142ppw@$      sq ~#y~�Aq ~ q ~1Et 143ppw@$      sq ~#y~�q ~ q ~1Et 144ppw@$      sq ~#y~��q ~ q ~1Et 145ppw@$      sq ~#y~�q ~ q ~1Et 146ppw@$      sq ~#y~�Eq ~ q ~1Et 147ppw@)v� �sq ~#y~�q ~ q ~1Et 148ppw@$      sq ~#y~��q ~ q ~1Et 149ppw@$      sq ~#y{_ �q ~ q ~1Et 15ppw@$      sq ~#y~?]q ~ q ~1Et 150ppw@$      sq ~#y~Cq ~ q ~1Et 151ppw@$      sq ~#y~F�q ~ q ~1Et 152ppw@(1���ssq ~#y~J�q ~ q ~1Et 153ppw@$      sq ~#y~Naq ~ q ~1Et 154ppw@*��&6�sq ~#y~R"q ~ q ~1Et 155ppw@$      sq ~#y~U�q ~ q ~1Et 156ppw@$      sq ~#y~Y�q ~ q ~1Et 157ppw@$      sq ~#y~]eq ~ q ~1Et 158ppw@$      sq ~#y~a&q ~ q ~1Et 159ppw@$      sq ~#y{_�q ~ q ~1Et 16ppw@$      sq ~#y~��q ~ q ~1Et 160ppw@$      sq ~#y~�}q ~ q ~1Et 161ppw@-����ńsq ~#y~�>q ~ q ~1Et 162ppw@-����ŀsq ~#y~��q ~ q ~1Et 163ppw@$      sq ~#y~��q ~ q ~1Et 164ppw@$      sq ~#y~Ɓq ~ q ~1Et 165ppw@%��9�}qsq ~#y~�Bq ~ q ~1Et 166ppw@$      sq ~#y~�q ~ q ~1Et 167ppw@&eNO���sq ~#y~��q ~ q ~1Et 168ppw@&Q�0��sq ~#y~Յq ~ q ~1Et 169ppw@$      sq ~#y{_wq ~ q ~1Et 17ppw@$      sq ~#y~(q ~ q ~1Et 170ppw@$      sq ~#y~+�q ~ q ~1Et 171ppw@$      sq ~#y~/�q ~ q ~1Et 172ppw@$      sq ~#y~3^q ~ q ~1Et 173ppw@$      sq ~#y~7q ~ q ~1Et 174ppw@$      sq ~#y~:�q ~ q ~1Et 175ppw@���h_�sq ~#y~>�q ~ q ~1Et 176ppw@$      sq ~#y~Bbq ~ q ~1Et 177ppw@$      sq ~#y~F#q ~ q ~1Et 178ppw@$      sq ~#y~I�q ~ q ~1Et 179ppw@$      sq ~#y{_8q ~ q ~1Et 18ppw@$      sq ~#y~�zq ~ q ~1Et 180ppw@$      sq ~#y~�;q ~ q ~1Et 181ppw@$      sq ~#y~��q ~ q ~1Et 182ppw@$      sq ~#y~��q ~ q ~1Et 183ppw@$      sq ~#y~�~q ~ q ~1Et 184ppw@$      sq ~#y~�?q ~ q ~1Et 185ppw@$      sq ~#y~� q ~ q ~1Et 186ppw@$      sq ~#y~��q ~ q ~1Et 187ppw@$      sq ~#y~��q ~ q ~1Et 188ppw@$      sq ~#y~�Cq ~ q ~1Et 189ppw@$      sq ~#y{_�q ~ q ~1Et 19ppw@%��9�}qsq ~#y~�q ~ q ~1Et 190ppw@5v��n�sq ~#y~�q ~ q ~1Et 191ppw@$      sq ~#y~[q ~ q ~1Et 192ppw@$      sq ~#y~q ~ q ~1Et 193ppw@$      sq ~#y~�q ~ q ~1Et 194ppw@$      sq ~#y~#�q ~ q ~1Et 195ppw@$      sq ~#y~'_q ~ q ~1Et 196ppw@$      sq ~#y~+ q ~ q ~1Et 197ppw@$      sq ~#y~.�q ~ q ~1Et 198ppw@$      sq ~#y~2�q ~ q ~1Et 199ppw@$      sq ~#y{H��q ~ q ~1Et 2ppw@$      sq ~#y{_b�q ~ q ~1Et 20ppw@$      sq ~#y~q ~ q ~1Et 200ppw@$      sq ~#y~�q ~ q ~1Et 201ppw@$      sq ~#y~�q ~ q ~1Et 202ppw@$      sq ~#y~Fq ~ q ~1Et 203ppw@$      sq ~#y~ q ~ q ~1Et 204ppw@'���@nsq ~#y~#�q ~ q ~1Et 205ppw@$      sq ~#y~'�q ~ q ~1Et 206ppw@$      sq ~#y~+Jq ~ q ~1Et 207ppw@$      sq ~#y~/q ~ q ~1Et 208ppw@$      sq ~#y~2�q ~ q ~1Et 209ppw@$      sq ~#y{_fPq ~ q ~1Et 21ppw@$      sq ~#y~�bq ~ q ~1Et 210ppw@$      sq ~#y~�#q ~ q ~1Et 211ppw@$      sq ~#y~��q ~ q ~1Et 212ppw@$      sq ~#y~��q ~ q ~1Et 213ppw@$      sq ~#y~�fq ~ q ~1Et 214ppw@$      sq ~#y~�'q ~ q ~1Et 215ppw@$      sq ~#y~��q ~ q ~1Et 216ppw@$      sq ~#y~��q ~ q ~1Et 217ppw@$      sq ~#y~�jq ~ q ~1Et 218ppw@$      sq ~#y~�+q ~ q ~1Et 219ppw@$      sq ~#y{_jq ~ q ~1Et 22ppw@$      sq ~#y~��q ~ q ~1Et 220ppw@$      sq ~#y~��q ~ q ~1Et 221ppw@$      sq ~#y~ Cq ~ q ~1Et 222ppw@$      sq ~#y~ q ~ q ~1Et 223ppw@$      sq ~#y~ �q ~ q ~1Et 224ppw@$      sq ~#y~ �q ~ q ~1Et 225ppw@$      sq ~#y~ Gq ~ q ~1Et 226ppw@$      sq ~#y~ q ~ q ~1Et 227ppw@$      sq ~#y~ �q ~ q ~1Et 228ppw@%Sx�d��sq ~#y~ �q ~ q ~1Et 229ppw@$      sq ~#y{_m�q ~ q ~1Et 23ppw@$      sq ~#y~ n q ~ q ~1Et 230ppw@$      sq ~#y~ q�q ~ q ~1Et 231ppw@$      sq ~#y~ u�q ~ q ~1Et 232ppw@$      sq ~#y~ ycq ~ q ~1Et 233ppw@$      sq ~#y~ }$q ~ q ~1Et 234ppw@$      sq ~#y~ ��q ~ q ~1Et 235ppw@$      sq ~#y~ ��q ~ q ~1Et 236ppw@$      sq ~#y~ �gq ~ q ~1Et 237ppw@$      sq ~#y~ �(q ~ q ~1Et 238ppw@$      sq ~#y~ ��q ~ q ~1Et 239ppw@$      sq ~#y{_q�q ~ q ~1Et 24ppw@$      sq ~#y~ �q ~ q ~1Et 240ppw@$      sq ~#y~ �@q ~ q ~1Et 241ppw@$      sq ~#y~ �q ~ q ~1Et 242ppw@$      sq ~#y~ ��q ~ q ~1Et 243ppw@$      sq ~#y~ �q ~ q ~1Et 244ppw@$      sq ~#y~ �Dq ~ q ~1Et 245ppw@$      sq ~#y~ �q ~ q ~1Et 246ppw@$      sq ~#y~ ��q ~ q ~1Et 247ppw@%U�e�W�sq ~#y~! �q ~ q ~1Et 248ppw@$      sq ~#y~!Hq ~ q ~1Et 249ppw@$      sq ~#y{_uTq ~ q ~1Et 25ppw@$      sq ~#y~!V�q ~ q ~1Et 250ppw@$      sq ~#y~!Z�q ~ q ~1Et 251ppw@$      sq ~#y~!^`q ~ q ~1Et 252ppw@$      sq ~#y~!b!q ~ q ~1Et 253ppw@$      sq ~#y~!e�q ~ q ~1Et 254ppw@5G�(��sq ~#y~!i�q ~ q ~1Et 255ppw@$      sq ~#y~!mdq ~ q ~1Et 256ppw@$      sq ~#y~!q%q ~ q ~1Et 257ppw@$      sq ~#y~!t�q ~ q ~1Et 258ppw@$      sq ~#y~!x�q ~ q ~1Et 259ppw@$      sq ~#y{_yq ~ q ~1Et 26ppw@$      sq ~#y~!�=q ~ q ~1Et 260ppw@ �Q,4�sq ~#y~!��q ~ q ~1Et 261ppw@$      sq ~#y~!ҿq ~ q ~1Et 262ppw@i���sq ~#y~!րq ~ q ~1Et 263ppw@$      sq ~#y~!�Aq ~ q ~1Et 264ppw@$      sq ~#y~!�q ~ q ~1Et 265ppw@$      sq ~#y~!��q ~ q ~1Et 266ppw@$      sq ~#y~!�q ~ q ~1Et 267ppw@$      sq ~#y~!�Eq ~ q ~1Et 268ppw@$      sq ~#y~!�q ~ q ~1Et 269ppw@$      sq ~#y{_|�q ~ q ~1Et 27ppw@$o� �@�sq ~#y~"?�q ~ q ~1Et 270ppw@$      sq ~#y~"C]q ~ q ~1Et 271ppw@$      sq ~#y~"Gq ~ q ~1Et 272ppw@@{5c�sq ~#y~"J�q ~ q ~1Et 273ppw@$      sq ~#y~"N�q ~ q ~1Et 274ppw@$      sq ~#y~"Raq ~ q ~1Et 275ppw@$      sq ~#y~"V"q ~ q ~1Et 276ppw@$      sq ~#y~"Y�q ~ q ~1Et 277ppw@$      sq ~#y~"]�q ~ q ~1Et 278ppw@$      sq ~#y~"aeq ~ q ~1Et 279ppw@$      sq ~#y{_��q ~ q ~1Et 28ppw@$      sq ~#y~"��q ~ q ~1Et 280ppw@$      sq ~#y~"��q ~ q ~1Et 281ppw@$      sq ~#y~"�}q ~ q ~1Et 282ppw@$      sq ~#y~"�>q ~ q ~1Et 283ppw@$      sq ~#y~"��q ~ q ~1Et 284ppw@$      sq ~#y~"��q ~ q ~1Et 285ppw@$      sq ~#y~"ʁq ~ q ~1Et 286ppw@$      sq ~#y~"�Bq ~ q ~1Et 287ppw@$      sq ~#y~"�q ~ q ~1Et 288ppw@$      sq ~#y~"��q ~ q ~1Et 289ppw@$      sq ~#y{_�Xq ~ q ~1Et 29ppw@$      sq ~#y~#(Zq ~ q ~1Et 290ppw@$      sq ~#y~#,q ~ q ~1Et 291ppw@$      sq ~#y~#/�q ~ q ~1Et 292ppw@$      sq ~#y~#3�q ~ q ~1Et 293ppw@$      sq ~#y~#7^q ~ q ~1Et 294ppw@$      sq ~#y~#;q ~ q ~1Et 295ppw@$      sq ~#y~#>�q ~ q ~1Et 296ppw@$      sq ~#y~#B�q ~ q ~1Et 297ppw@$      sq ~#y~#Fbq ~ q ~1Et 298ppw@$      sq ~#y~#J#q ~ q ~1Et 299ppw@$      sq ~#y{H�Dq ~ q ~1Et 3ppw@$      sq ~#y{_��q ~ q ~1Et 30ppw@$      sq ~#y~-(�q ~ q ~1Et 300ppw@$      sq ~#y~-,Eq ~ q ~1Et 301ppw@$      sq ~#y~-0q ~ q ~1Et 302ppw@$      sq ~#y~-3�q ~ q ~1Et 303ppw@$      sq ~#y~-7�q ~ q ~1Et 304ppw@$      sq ~#y~-;Iq ~ q ~1Et 305ppw@$      sq ~#y~-?
q ~ q ~1Et 306ppw@$      sq ~#y~-B�q ~ q ~1Et 307ppw@$      sq ~#y~-F�q ~ q ~1Et 308ppw@$      sq ~#y~-JMq ~ q ~1Et 309ppw@$      sq ~#y{_گq ~ q ~1Et 31ppw@$      sq ~#y~-��q ~ q ~1Et 310ppw@$      sq ~#y~-��q ~ q ~1Et 311ppw@$      sq ~#y~-�eq ~ q ~1Et 312ppw@$      sq ~#y~-�&q ~ q ~1Et 313ppw@$      sq ~#y~-��q ~ q ~1Et 314ppw@$      sq ~#y~-��q ~ q ~1Et 315ppw@$      sq ~#y~-�iq ~ q ~1Et 316ppw@$      sq ~#y~-�*q ~ q ~1Et 317ppw@$      sq ~#y~-��q ~ q ~1Et 318ppw@$      sq ~#y~-��q ~ q ~1Et 319ppw@$      sq ~#y{_�pq ~ q ~1Et 32ppw@$      sq ~#y~.Bq ~ q ~1Et 320ppw@$      sq ~#y~.q ~ q ~1Et 321ppw@$      sq ~#y~.�q ~ q ~1Et 322ppw@$      sq ~#y~.�q ~ q ~1Et 323ppw@$      sq ~#y~. Fq ~ q ~1Et 324ppw@$      sq ~#y~.$q ~ q ~1Et 325ppw@$      sq ~#y~.'�q ~ q ~1Et 326ppw@$      sq ~#y~.+�q ~ q ~1Et 327ppw@$      sq ~#y~./Jq ~ q ~1Et 328ppw@$      sq ~#y~.3q ~ q ~1Et 329ppw@$      sq ~#y{_�1q ~ q ~1Et 33ppw@$      sq ~#y~.��q ~ q ~1Et 330ppw@$      sq ~#y~.�bq ~ q ~1Et 331ppw@$      sq ~#y~.�#q ~ q ~1Et 332ppw@$      sq ~#y~.��q ~ q ~1Et 333ppw@$      sq ~#y~.��q ~ q ~1Et 334ppw@$      sq ~#y~.�fq ~ q ~1Et 335ppw@$      sq ~#y~.�'q ~ q ~1Et 336ppw@$      sq ~#y~.��q ~ q ~1Et 337ppw@$      sq ~#y~.��q ~ q ~1Et 338ppw@$      sq ~#y~.�jq ~ q ~1Et 339ppw@$      sq ~#y{_��q ~ q ~1Et 34ppw@$      sq ~#y~.� q ~ q ~1Et 340ppw@$      sq ~#y~.��q ~ q ~1Et 341ppw@$      sq ~#y~/�q ~ q ~1Et 342ppw@$      sq ~#y~/Cq ~ q ~1Et 343ppw@$      sq ~#y~/	q ~ q ~1Et 344ppw@$      sq ~#y~/�q ~ q ~1Et 345ppw@i���sq ~#y~/�q ~ q ~1Et 346ppw@$      sq ~#y~/Gq ~ q ~1Et 347ppw@$      sq ~#y~/q ~ q ~1Et 348ppw@$      sq ~#y~/�q ~ q ~1Et 349ppw@$      sq ~#y{_�q ~ q ~1Et 35ppw@$      sq ~#y~/n_q ~ q ~1Et 350ppw@-����ŀsq ~#y~/r q ~ q ~1Et 351ppw@$      sq ~#y~/u�q ~ q ~1Et 352ppw@$      sq ~#y~/y�q ~ q ~1Et 353ppw@$      sq ~#y~/}cq ~ q ~1Et 354ppw@$      sq ~#y~/�$q ~ q ~1Et 355ppw@$      sq ~#y~/��q ~ q ~1Et 356ppw@$      sq ~#y~/��q ~ q ~1Et 357ppw@$      sq ~#y~/�gq ~ q ~1Et 358ppw@$      sq ~#y~/�(q ~ q ~1Et 359ppw@$      sq ~#y{_�tq ~ q ~1Et 36ppw@$      sq ~#y~/�q ~ q ~1Et 360ppw@$      sq ~#y~/�q ~ q ~1Et 361ppw@$      sq ~#y~/�@q ~ q ~1Et 362ppw@$      sq ~#y~/�q ~ q ~1Et 363ppw@$      sq ~#y~/��q ~ q ~1Et 364ppw@ �̾�,sq ~#y~/��q ~ q ~1Et 365ppw@$      sq ~#y~/�Dq ~ q ~1Et 366ppw@$      sq ~#y~/�q ~ q ~1Et 367ppw@$      sq ~#y~0 �q ~ q ~1Et 368ppw@$      sq ~#y~0�q ~ q ~1Et 369ppw@%��9�}qsq ~#y{_�5q ~ q ~1Et 37ppw@#��吢sq ~#y~0Wq ~ q ~1Et 370ppw@$      sq ~#y~0Z�q ~ q ~1Et 371ppw@$      sq ~#y~0^�q ~ q ~1Et 372ppw@$      sq ~#y~0b`q ~ q ~1Et 373ppw@&'��5V�sq ~#y~0f!q ~ q ~1Et 374ppw@$      sq ~#y~0i�q ~ q ~1Et 375ppw@$      sq ~#y~0m�q ~ q ~1Et 376ppw@$      sq ~#y~0qdq ~ q ~1Et 377ppw@$      sq ~#y~0u%q ~ q ~1Et 378ppw@$      sq ~#y~0x�q ~ q ~1Et 379ppw@$      sq ~#y{_��q ~ q ~1Et 38ppw@$      sq ~#y~0�|q ~ q ~1Et 380ppw@$      sq ~#y~0�=q ~ q ~1Et 381ppw@$      sq ~#y~0��q ~ q ~1Et 382ppw@$      sq ~#y~0ֿq ~ q ~1Et 383ppw@$      sq ~#y~0ڀq ~ q ~1Et 384ppw@$      sq ~#y~0�Aq ~ q ~1Et 385ppw@$      sq ~#y~0�q ~ q ~1Et 386ppw@$      sq ~#y~0��q ~ q ~1Et 387ppw@$      sq ~#y~0�q ~ q ~1Et 388ppw@$      sq ~#y~0�Eq ~ q ~1Et 389ppw@$      sq ~#y{_��q ~ q ~1Et 39ppw@$      sq ~#y~1?�q ~ q ~1Et 390ppw@$      sq ~#y~1C�q ~ q ~1Et 391ppw@$      sq ~#y~1G]q ~ q ~1Et 392ppw@$      sq ~#y~1Kq ~ q ~1Et 393ppw@$      sq ~#y~1N�q ~ q ~1Et 394ppw@$      sq ~#y~1R�q ~ q ~1Et 395ppw@$      sq ~#y~1Vaq ~ q ~1Et 396ppw@$      sq ~#y~1Z"q ~ q ~1Et 397ppw@$      sq ~#y~1]�q ~ q ~1Et 398ppw@$      sq ~#y~1a�q ~ q ~1Et 399ppw@$      sq ~#y{H�q ~ q ~1Et 4ppw@(L*�c�sq ~#y{`KMq ~ q ~1Et 40ppw@5v��n�sq ~#y~;@q ~ q ~1Et 400ppw@$      sq ~#y~;C�q ~ q ~1Et 401ppw@$      sq ~#y~;G�q ~ q ~1Et 402ppw@$      sq ~#y~;KHq ~ q ~1Et 403ppw@$      sq ~#y~;O	q ~ q ~1Et 404ppw@$      sq ~#y~;R�q ~ q ~1Et 405ppw@$      sq ~#y~;V�q ~ q ~1Et 406ppw@$      sq ~#y~;ZLq ~ q ~1Et 407ppw@$      sq ~#y~;^q ~ q ~1Et 408ppw@$      sq ~#y~;a�q ~ q ~1Et 409ppw@$      sq ~#y{`Oq ~ q ~1Et 41ppw@$      sq ~#y~;�dq ~ q ~1Et 410ppw@$      sq ~#y~;�%q ~ q ~1Et 411ppw@$      sq ~#y~;��q ~ q ~1Et 412ppw@$      sq ~#y~;��q ~ q ~1Et 413ppw@$      sq ~#y~;�hq ~ q ~1Et 414ppw@$      sq ~#y~;�)q ~ q ~1Et 415ppw@$      sq ~#y~;��q ~ q ~1Et 416ppw@$      sq ~#y~;Ϋq ~ q ~1Et 417ppw@$      sq ~#y~;�lq ~ q ~1Et 418ppw@$      sq ~#y~;�-q ~ q ~1Et 419ppw@$      sq ~#y{`R�q ~ q ~1Et 42ppw@$      sq ~#y~<(�q ~ q ~1Et 420ppw@$      sq ~#y~<,�q ~ q ~1Et 421ppw@$      sq ~#y~<0Eq ~ q ~1Et 422ppw@$      sq ~#y~<4q ~ q ~1Et 423ppw@$      sq ~#y~<7�q ~ q ~1Et 424ppw@$      sq ~#y~<;�q ~ q ~1Et 425ppw@$      sq ~#y~<?Iq ~ q ~1Et 426ppw@$      sq ~#y~<C
q ~ q ~1Et 427ppw@$      sq ~#y~<F�q ~ q ~1Et 428ppw@$      sq ~#y~<J�q ~ q ~1Et 429ppw@�iu��sq ~#y{`V�q ~ q ~1Et 43ppw@$�g\oQsq ~#y~<�"q ~ q ~1Et 430ppw@$����sq ~#y~<��q ~ q ~1Et 431ppw?��2Q�v�sq ~#y~<��q ~ q ~1Et 432ppw@�xJdGsq ~#y~<�eq ~ q ~1Et 433ppw@$��D��asq ~#y~<�&q ~ q ~1Et 434ppw@�<�hG�sq ~#y~<��q ~ q ~1Et 435ppw?��s��֓sq ~#y~<��q ~ q ~1Et 436ppw?��s��֓sq ~#y~<�iq ~ q ~1Et 437ppw@sw�:sq ~#y~<�*q ~ q ~1Et 438ppw@���Nsq ~#y{`ZQq ~ q ~1Et 44ppw@$      sq ~#y{`^q ~ q ~1Et 45ppw@$      sq ~#y{`a�q ~ q ~1Et 46ppw@$      sq ~#y{`e�q ~ q ~1Et 47ppw@$      sq ~#y{`iUq ~ q ~1Et 48ppw@$�g\oIsq ~#y{`mq ~ q ~1Et 49ppw@$      sq ~#y{H��q ~ q ~1Et 5ppw@$      sq ~#y{`��q ~ q ~1Et 50ppw@$      sq ~#y{`�mq ~ q ~1Et 51ppw@$      sq ~#y{`�.q ~ q ~1Et 52ppw@$      sq ~#y{`��q ~ q ~1Et 53ppw@$      sq ~#y{`ΰq ~ q ~1Et 54ppw@$      sq ~#y{`�qq ~ q ~1Et 55ppw@$      sq ~#y{`�2q ~ q ~1Et 56ppw@$      sq ~#y{`��q ~ q ~1Et 57ppw@$      sq ~#y{`ݴq ~ q ~1Et 58ppw@$      sq ~#y{`�uq ~ q ~1Et 59ppw@���h_�sq ~#y{H��q ~ q ~1Et 6ppw@$      sq ~#y{a4q ~ q ~1Et 60ppw@���h_�sq ~#y{a7�q ~ q ~1Et 61ppw@$      sq ~#y{a;�q ~ q ~1Et 62ppw@$      sq ~#y{a?Nq ~ q ~1Et 63ppw@$      sq ~#y{aCq ~ q ~1Et 64ppw@$      sq ~#y{aF�q ~ q ~1Et 65ppw@$      sq ~#y{aJ�q ~ q ~1Et 66ppw@$      sq ~#y{aNRq ~ q ~1Et 67ppw@$      sq ~#y{aRq ~ q ~1Et 68ppw@$      sq ~#y{aU�q ~ q ~1Et 69ppw@#�
2!�sq ~#y{H�Hq ~ q ~1Et 7ppw@$      sq ~#y{a�jq ~ q ~1Et 70ppw@$      sq ~#y{a�+q ~ q ~1Et 71ppw@$      sq ~#y{a��q ~ q ~1Et 72ppw@$      sq ~#y{a��q ~ q ~1Et 73ppw@$      sq ~#y{a�nq ~ q ~1Et 74ppw@$      sq ~#y{a�/q ~ q ~1Et 75ppw@$      sq ~#y{a��q ~ q ~1Et 76ppw@$      sq ~#y{a±q ~ q ~1Et 77ppw@$      sq ~#y{a�rq ~ q ~1Et 78ppw@$      sq ~#y{a�3q ~ q ~1Et 79ppw@$      sq ~#y{H�	q ~ q ~1Et 8ppw@$      sq ~#y{b�q ~ q ~1Et 80ppw@$      sq ~#y{b �q ~ q ~1Et 81ppw@$      sq ~#y{b$Kq ~ q ~1Et 82ppw@$      sq ~#y{b(q ~ q ~1Et 83ppw@$      sq ~#y{b+�q ~ q ~1Et 84ppw@$      sq ~#y{b/�q ~ q ~1Et 85ppw@$      sq ~#y{b3Oq ~ q ~1Et 86ppw@$      sq ~#y{b7q ~ q ~1Et 87ppw@$      sq ~#y{b:�q ~ q ~1Et 88ppw@$      sq ~#y{b>�q ~ q ~1Et 89ppw@$      sq ~#y{H��q ~ q ~1Et 9ppw@$      sq ~#y{b�(q ~ q ~1Et 90ppw@$      sq ~#y{b��q ~ q ~1Et 91ppw@$      sq ~#y{b��q ~ q ~1Et 92ppw@$      sq ~#y{b�kq ~ q ~1Et 93ppw@$      sq ~#y{b�,q ~ q ~1Et 94ppw@$      sq ~#y{b��q ~ q ~1Et 95ppw@$      sq ~#y{b��q ~ q ~1Et 96ppw@$      sq ~#y{b�oq ~ q ~1Et 97ppw@$      sq ~#y{b�0q ~ q ~1Et 98ppw@i���sq ~#y{b��q ~ q ~1Et 99ppw@$      q ~#|w?�      sq ~#y��u�t LOGEXPt CPP1q ~Oq ~nq ~ Dw@QS}�sq ~#yd!+�t RULEt <applypppw?���bP��sq ~#y��	�q ~4�t >applypppw@�ܓk*Qsq ~#y4::�q ~4�t 	>thatlesspppw?�g�-�hsq ~#yZ�q ~4�t >trcomp1pppw?��C,� �sq ~#yԿq ~4�t lexpppw@#�-��sq ~#yR롞q ~4�t shift_pppppw��i�n]�x